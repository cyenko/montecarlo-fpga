----------------------------------------------------------------------------- 
library IEEE; 
 
use IEEE.std_logic_1164.all; 
use WORK.monte_carlo.all; 
--Additional standard or custom libraries go here 
use IEEE.numeric_std.all;

--inputs: clock, start, stock price, strike, t
--output: premium, stock price out, ready
--	for now, do only premium and ready

entity sqrt_fn is 
 port( 
	 --Inputs (is unsigned)
	 clk : in std_logic; 
	 bitVector : in std_logic_vector (7 downto 0); --8 bits
	 
	 --Outputs (is fixed point)
	 outVector : out std_logic_vector (15 downto 0)
 ); 
end entity sqrt_fn;

architecture behavioral of sqrt_fn is 
--Declare the ROM type
--Real length will be 0 to 2**16-1
--type rom is array (0 to (2**16)-1) of std_logic_vector(15 downto 0);
type rom is array (0 to (127)) of std_logic_vector(15 downto 0);
--Input the LUT, this will be generated by python
constant sqrt_lut : rom := (0 => "0000000000000000",
1 => "0000000100000000",2 => "0000000101101010",3 => "0000000110111011",
4 => "0000001000000000",5 => "0000001000111100",6 => "0000001001110011",
7 => "0000001010100101",8 => "0000001011010100",9 => "0000001100000000",
10 => "0000001100101001",11 => "0000001101010001",12 => "0000001101110110",
13 => "0000001110011011",14 => "0000001110111101",15 => "0000001111011111",
16 => "0000010000000000",17 => "0000010000011111",18 => "0000010000111110",
19 => "0000010001011011",20 => "0000010001111000",21 => "0000010010010101",
22 => "0000010010110000",23 => "0000010011001011",24 => "0000010011100110",
25 => "0000010100000000",26 => "0000010100011001",27 => "0000010100110010",
28 => "0000010101001010",29 => "0000010101100010",30 => "0000010101111010",
31 => "0000010110010001",32 => "0000010110101000",33 => "0000010110111110",
34 => "0000010111010100",35 => "0000010111101010",36 => "0000011000000000",
37 => "0000011000010101",38 => "0000011000101010",39 => "0000011000111110",
40 => "0000011001010011",41 => "0000011001100111",42 => "0000011001111011",
43 => "0000011010001110",44 => "0000011010100010",45 => "0000011010110101",
46 => "0000011011001000",47 => "0000011011011011",48 => "0000011011101101",
49 => "0000011100000000",50 => "0000011100010010",51 => "0000011100100100",
52 => "0000011100110110",53 => "0000011101000111",54 => "0000011101011001",
55 => "0000011101101010",56 => "0000011101111011",57 => "0000011110001100",
58 => "0000011110011101",59 => "0000011110101110",60 => "0000011110111110",
61 => "0000011111001111",62 => "0000011111011111",63 => "0000011111101111",
64 => "0000100000000000",65 => "0000100000001111",66 => "0000100000011111",
67 => "0000100000101111",68 => "0000100000111111",69 => "0000100001001110",
70 => "0000100001011101",71 => "0000100001101101",72 => "0000100001111100",
73 => "0000100010001011",74 => "0000100010011010",75 => "0000100010101001",
76 => "0000100010110111",77 => "0000100011000110",78 => "0000100011010100",
79 => "0000100011100011",80 => "0000100011110001",81 => "0000100100000000",
82 => "0000100100001110",83 => "0000100100011100",84 => "0000100100101010",
85 => "0000100100111000",86 => "0000100101000110",87 => "0000100101010011",
88 => "0000100101100001",89 => "0000100101101111",90 => "0000100101111100",
91 => "0000100110001010",92 => "0000100110010111",93 => "0000100110100100",
94 => "0000100110110010",95 => "0000100110111111",96 => "0000100111001100",
97 => "0000100111011001",98 => "0000100111100110",99 => "0000100111110011",
100 => "0000101000000000",101 => "0000101000001100",102 => "0000101000011001",
103 => "0000101000100110",104 => "0000101000110010",105 => "0000101000111111",
106 => "0000101001001011",107 => "0000101001011000",108 => "0000101001100100",
109 => "0000101001110000",110 => "0000101001111100",111 => "0000101010001001",
112 => "0000101010010101",113 => "0000101010100001",114 => "0000101010101101",
115 => "0000101010111001",116 => "0000101011000101",117 => "0000101011010001",
118 => "0000101011011100",119 => "0000101011101000",120 => "0000101011110100",
121 => "0000101100000000",122 => "0000101100001011",123 => "0000101100010111",
124 => "0000101100100010",125 => "0000101100101110",126 => "0000101100111001",
127 => "0000101101000100");

begin

	findValue: process (clk,bitVector) is 
		variable index : integer := 0;

		BEGIN  
			index := to_integer(unsigned(bitVector));
			if index < 127 then
				outVector <= sqrt_lut(index);
			else 
				outVector <= x"0000";
			end if;

	end process findValue;

end architecture;

