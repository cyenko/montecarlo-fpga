----------------------------------------------------------------------------- 
library IEEE; 
 
use IEEE.std_logic_1164.all; 
use WORK.monte_carlo.all; 
--Additional standard or custom libraries go here 
use IEEE.numeric_std.all;

--inputs: clock, start, stock price, strike, t
--output: premium, stock price out, ready
--	for now, do only premium and ready

entity exp is 
 port( 
	 --Inputs 
	 clk : in std_logic; 
	 bitVector : in std_logic_vector (15 downto 0); --16 bits
	 
	 --Outputs 
	 outVector : out std_logic_vector (15 downto 0)
 ); 
end entity exp;

architecture behavioral of exp is 
--Declare the ROM type
--Real length will be 0 to 2**16-1
type rom is array (0 to (2**16)-1) of std_logic_vector(15 downto 0);
--Input the LUT, this will be generated by python
--constant exp_lut : rom := (0=>"0000000000000000",1=>"0000000000000001");
constant exp_lut : rom := (0 => "0000100000000000",
1 => "0000100001101001",2 => "0000100011011101",
3 => "0000100000100011",4 => "0000100111101100",
5 => "0000101010001001",6 => "0000101100110110",
7 => "0001000000001110",8 => "0001000011100010",
9 => "0001000000101110",10 => "0000100001101001",
11 => "0000100001110100",12 => "0000100001111111",
13 => "0000100010001011",14 => "0000100000001111",
15 => "0000100010100010",16 => "0000100010101110",
17 => "0000100010111001",18 => "0000100011000101",
19 => "0000100011010001",20 => "0000100011011101",
21 => "0000100011101010",22 => "0000100011110110",
23 => "0000100100000011",24 => "0000100100001111",
25 => "0000100100011100",26 => "0000100100101001",
27 => "0000100000011111",28 => "0000100101000011",
29 => "0000100101010000",30 => "0000100000100011",
31 => "0000100101101011",32 => "0000100101111001",
33 => "0000100110000111",34 => "0000100110010101",
35 => "0000100110100011",36 => "0000100110110001",
37 => "0000100111000000",38 => "0000100111001110",
39 => "0000100111011101",40 => "0000100111101100",
41 => "0000100111111011",42 => "0000101000001010",
43 => "0000101000011001",44 => "0000101000101001",
45 => "0000101000111000",46 => "0000101001001000",
47 => "0000100000000110",48 => "0000101001101000",
49 => "0000101001111000",50 => "0000101010001001",
51 => "0000101010011001",52 => "0000101010101010",
53 => "0000101010111011",54 => "0000101011001100",
55 => "0000101011011101",56 => "0000101011101111",
57 => "0000101100000000",58 => "0000101100010010",
59 => "0000101100100100",60 => "0000101100110110",
61 => "0000100001010100",62 => "0000101101011011",
63 => "0000101101101110",64 => "0000101110000000",
65 => "0000101110010100",66 => "0000101110100111",
67 => "0000101110111010",68 => "0000101111001110",
69 => "0000101111100010",70 => "0001000000001110",
71 => "0001000000100010",72 => "0001000000110110",
73 => "0001000001001011",74 => "0001000001100000",
75 => "0001000001110101",76 => "0001000010001010",
77 => "0001000000010000",78 => "0001000010110101",
79 => "0001000011001011",80 => "0001000011100010",
81 => "0001000011111000",82 => "0001000000011011",
83 => "0001000100100101",84 => "0001000100111100",
85 => "0001000000100010",86 => "0001000101101011",
87 => "0001000110000011",88 => "0001000110011011",
89 => "0001000110110011",90 => "0001000000101110",
91 => "0001000111100100",92 => "0001000111111101",
93 => "0001001000010111",94 => "0001000000111000",
95 => "0001001001001010",96 => "0001001001100100",
97 => "0001001001111110",98 => "0001001010011000",
99 => "0001001010110011",100 => "0000100001101001",
101 => "0000100001101010",102 => "0000100001101011",
103 => "0000100001101100",104 => "0000100000001011",
105 => "0000100001101111",106 => "0000100001110000",
107 => "0000100001110001",108 => "0000100001110010",
109 => "0000100001110011",110 => "0000100001110100",
111 => "0000100001110101",112 => "0000100001110111",
113 => "0000100000001100",114 => "0000100001111001",
115 => "0000100001111010",116 => "0000100001111011",
117 => "0000100001111100",118 => "0000100001111101",
119 => "0000100001111110",120 => "0000100001111111",
121 => "0000100010000001",122 => "0000100000001101",
123 => "0000100010000011",124 => "0000100010000100",
125 => "0000100010000101",126 => "0000100010000110",
127 => "0000100010000111",128 => "0000100010001001",
129 => "0000100010001010",130 => "0000100010001011",
131 => "0000100000001110",132 => "0000100010001101",
133 => "0000100010001110",134 => "0000100010001111",
135 => "0000100010010001",136 => "0000100010010010",
137 => "0000100010010011",138 => "0000100010010100",
139 => "0000100010010101",140 => "0000100000001111",
141 => "0000100010010111",142 => "0000100010011001",
143 => "0000100010011010",144 => "0000100010011011",
145 => "0000100010011100",146 => "0000100010011101",
147 => "0000100010011110",148 => "0000100000010000",
149 => "0000100010100001",150 => "0000100010100010",
151 => "0000100010100011",152 => "0000100010100100",
153 => "0000100010100101",154 => "0000100010100110",
155 => "0000100010101000",156 => "0000100010101001",
157 => "0000100000010001",158 => "0000100010101011",
159 => "0000100010101100",160 => "0000100010101110",
161 => "0000100010101111",162 => "0000100010110000",
163 => "0000100010110001",164 => "0000100010110010",
165 => "0000100010110011",166 => "0000100010110101",
167 => "0000100010110110",168 => "0000100010110111",
169 => "0000100010111000",170 => "0000100010111001",
171 => "0000100010111010",172 => "0000100010111100",
173 => "0000100010111101",174 => "0000100000010011",
175 => "0000100010111111",176 => "0000100011000000",
177 => "0000100011000010",178 => "0000100011000011",
179 => "0000100011000100",180 => "0000100011000101",
181 => "0000100011000110",182 => "0000100000000010",
183 => "0000100011001001",184 => "0000100011001010",
185 => "0000100011001011",186 => "0000100011001100",
187 => "0000100011001110",188 => "0000100011001111",
189 => "0000100011010000",190 => "0000100011010001",
191 => "0000100000010101",192 => "0000100011010100",
193 => "0000100011010101",194 => "0000100011010110",
195 => "0000100011010111",196 => "0000100011011001",
197 => "0000100011011010",198 => "0000100011011011",
199 => "0000100000010110",200 => "0000100011011101",
201 => "0000100011011111",202 => "0000100011100000",
203 => "0000100011100001",204 => "0000100011100010",
205 => "0000100011100100",206 => "0000100011100101",
207 => "0000100000010111",208 => "0000100011100111",
209 => "0000100011101000",210 => "0000100011101010",
211 => "0000100011101011",212 => "0000100011101100",
213 => "0000100011101101",214 => "0000100011101111",
215 => "0000100000011000",216 => "0000100011110001",
217 => "0000100011110010",218 => "0000100011110100",
219 => "0000100011110101",220 => "0000100011110110",
221 => "0000100011110111",222 => "0000100011111001",
223 => "0000100000011001",224 => "0000100011111011",
225 => "0000100011111100",226 => "0000100011111110",
227 => "0000100011111111",228 => "0000100100000000",
229 => "0000100100000001",230 => "0000100100000011",
231 => "0000100000011010",232 => "0000100100000101",
233 => "0000100100000110",234 => "0000100100001000",
235 => "0000100100001001",236 => "0000100100001010",
237 => "0000100100001011",238 => "0000100100001101",
239 => "0000100000011011",240 => "0000100100001111",
241 => "0000100100010001",242 => "0000100100010010",
243 => "0000100100010011",244 => "0000100100010100",
245 => "0000100100010110",246 => "0000100100010111",
247 => "0000100000011100",248 => "0000100100011001",
249 => "0000100100011011",250 => "0000100100011100",
251 => "0000100100011101",252 => "0000100100011111",
253 => "0000100100100000",254 => "0000100100100001",
255 => "0000100000011101",256 => "0000100100100100",
257 => "0000100100100101",258 => "0000100100100110",
259 => "0000100100101000",260 => "0000100100101001",
261 => "0000100100101010",262 => "0000100000000011",
263 => "0000100100101101",264 => "0000100100101110",
265 => "0000100100101111",266 => "0000100100110001",
267 => "0000100100110010",268 => "0000100100110011",
269 => "0000100100110101",270 => "0000100000011111",
271 => "0000100100110111",272 => "0000100100111001",
273 => "0000100100111010",274 => "0000100100111011",
275 => "0000100100111101",276 => "0000100100111110",
277 => "0000100100111111",278 => "0000100000100000",
279 => "0000100101000010",280 => "0000100101000011",
281 => "0000100101000100",282 => "0000100101000110",
283 => "0000100101000111",284 => "0000100101001000",
285 => "0000100000100001",286 => "0000100101001011",
287 => "0000100101001100",288 => "0000100101001110",
289 => "0000100101001111",290 => "0000100101010000",
291 => "0000100101010010",292 => "0000100101010011",
293 => "0000100000100010",294 => "0000100101010110",
295 => "0000100101010111",296 => "0000100101011000",
297 => "0000100101011010",298 => "0000100101011011",
299 => "0000100101011101",300 => "0000100000100011",
301 => "0000100101011111",302 => "0000100101100001",
303 => "0000100101100010",304 => "0000100101100011",
305 => "0000100101100101",306 => "0000100101100110",
307 => "0000100101100111",308 => "0000100101101001",
309 => "0000100101101010",310 => "0000100101101011",
311 => "0000100101101101",312 => "0000100101101110",
313 => "0000100101110000",314 => "0000100101110001",
315 => "0000100000100101",316 => "0000100101110100",
317 => "0000100101110101",318 => "0000100101110110",
319 => "0000100101111000",320 => "0000100101111001",
321 => "0000100101111011",322 => "0000100000100110",
323 => "0000100101111101",324 => "0000100101111111",
325 => "0000100110000000",326 => "0000100110000001",
327 => "0000100110000011",328 => "0000100110000100",
329 => "0000100000100111",330 => "0000100110000111",
331 => "0000100110001000",332 => "0000100110001010",
333 => "0000100110001011",334 => "0000100110001101",
335 => "0000100110001110",336 => "0000100110001111",
337 => "0000100110010001",338 => "0000100110010010",
339 => "0000100110010100",340 => "0000100110010101",
341 => "0000100110010110",342 => "0000100110011000",
343 => "0000100110011001",344 => "0000100110011011",
345 => "0000100110011100",346 => "0000100110011101",
347 => "0000100110011111",348 => "0000100110100000",
349 => "0000100110100010",350 => "0000100110100011",
351 => "0000100000101010",352 => "0000100110100110",
353 => "0000100110100111",354 => "0000100110101001",
355 => "0000100110101010",356 => "0000100110101100",
357 => "0000100110101101",358 => "0000100000101011",
359 => "0000100110110000",360 => "0000100110110001",
361 => "0000100110110011",362 => "0000100110110100",
363 => "0000100110110110",364 => "0000100110110111",
365 => "0000100110111001",366 => "0000100110111010",
367 => "0000100110111011",368 => "0000100110111101",
369 => "0000100110111110",370 => "0000100111000000",
371 => "0000100111000001",372 => "0000100111000011",
373 => "0000100111000100",374 => "0000100111000110",
375 => "0000100111000111",376 => "0000100111001000",
377 => "0000100111001010",378 => "0000100111001011",
379 => "0000100111001101",380 => "0000100111001110",
381 => "0000100111010000",382 => "0000100111010001",
383 => "0000100111010011",384 => "0000100111010100",
385 => "0000100000101111",386 => "0000100111010111",
387 => "0000100111011001",388 => "0000100111011010",
389 => "0000100111011100",390 => "0000100111011101",
391 => "0000100111011110",392 => "0000100000110000",
393 => "0000100111100001",394 => "0000100111100011",
395 => "0000100111100100",396 => "0000100111100110",
397 => "0000100111100111",398 => "0000100111101001",
399 => "0000100000110001",400 => "0000100111101100",
401 => "0000100111101101",402 => "0000100111101111",
403 => "0000100111110000",404 => "0000100111110010",
405 => "0000100111110011",406 => "0000100111110101",
407 => "0000100111110110",408 => "0000100111111000",
409 => "0000100111111001",410 => "0000100111111011",
411 => "0000100111111100",412 => "0000100000110011",
413 => "0000100111111111",414 => "0000101000000001",
415 => "0000101000000010",416 => "0000101000000100",
417 => "0000101000000101",418 => "0000101000000111",
419 => "0000100000110100",420 => "0000101000001010",
421 => "0000101000001011",422 => "0000101000001101",
423 => "0000101000001111",424 => "0000101000010000",
425 => "0000100000110101",426 => "0000101000010011",
427 => "0000101000010101",428 => "0000101000010110",
429 => "0000101000011000",430 => "0000101000011001",
431 => "0000101000011011",432 => "0000100000110110",
433 => "0000101000011110",434 => "0000101000011111",
435 => "0000101000100001",436 => "0000101000100011",
437 => "0000101000100100",438 => "0000100000110111",
439 => "0000101000100111",440 => "0000101000101001",
441 => "0000101000101010",442 => "0000101000101100",
443 => "0000101000101101",444 => "0000101000101111",
445 => "0000100000111000",446 => "0000101000110010",
447 => "0000101000110100",448 => "0000101000110101",
449 => "0000101000110111",450 => "0000101000111000",
451 => "0000100000111001",452 => "0000101000111011",
453 => "0000101000111101",454 => "0000101000111111",
455 => "0000101001000000",456 => "0000101001000010",
457 => "0000101001000011",458 => "0000101001000101",
459 => "0000101001000110",460 => "0000101001001000",
461 => "0000101001001010",462 => "0000101001001011",
463 => "0000101001001101",464 => "0000100000111011",
465 => "0000101001010000",466 => "0000101001010010",
467 => "0000101001010011",468 => "0000101001010101",
469 => "0000101001010110",470 => "0000100000000110",
471 => "0000101001011010",472 => "0000101001011011",
473 => "0000101001011101",474 => "0000101001011110",
475 => "0000101001100000",476 => "0000100000111101",
477 => "0000101001100011",478 => "0000101001100101",
479 => "0000101001100110",480 => "0000101001101000",
481 => "0000101001101010",482 => "0000101001101011",
483 => "0000101001101101",484 => "0000101001101111",
485 => "0000101001110000",486 => "0000101001110010",
487 => "0000101001110011",488 => "0000101001110101",
489 => "0000101001110111",490 => "0000101001111000",
491 => "0000101001111010",492 => "0000101001111100",
493 => "0000101001111101",494 => "0000101001111111",
495 => "0000100001000000",496 => "0000101010000010",
497 => "0000101010000100",498 => "0000101010000101",
499 => "0000101010000111",500 => "0000101010001001",
501 => "0000100001000001",502 => "0000101010001100",
503 => "0000101010001110",504 => "0000101010001111",
505 => "0000101010010001",506 => "0000101010010011",
507 => "0000100001000010",508 => "0000101010010110",
509 => "0000101010011000",510 => "0000101010011001",
511 => "0000101010011011",512 => "0000101010011101",
513 => "0000100001000011",514 => "0000101010100000",
515 => "0000101010100010",516 => "0000101010100011",
517 => "0000101010100101",518 => "0000101010100111",
519 => "0000100001000100",520 => "0000101010101010",
521 => "0000101010101100",522 => "0000101010101101",
523 => "0000101010101111",524 => "0000101010110001",
525 => "0000100001000101",526 => "0000101010110100",
527 => "0000101010110110",528 => "0000101010111000",
529 => "0000101010111001",530 => "0000101010111011",
531 => "0000101010111101",532 => "0000101010111110",
533 => "0000101011000000",534 => "0000101011000010",
535 => "0000101011000011",536 => "0000101011000101",
537 => "0000101011000111",538 => "0000101011001001",
539 => "0000101011001010",540 => "0000101011001100",
541 => "0000101011001110",542 => "0000101011001111",
543 => "0000101011010001",544 => "0000101011010011",
545 => "0000101011010101",546 => "0000101011010110",
547 => "0000101011011000",548 => "0000100001001001",
549 => "0000101011011100",550 => "0000101011011101",
551 => "0000101011011111",552 => "0000101011100001",
553 => "0000101011100010",554 => "0000100001001010",
555 => "0000101011100110",556 => "0000101011101000",
557 => "0000101011101001",558 => "0000101011101011",
559 => "0000101011101101",560 => "0000101011101111",
561 => "0000101011110000",562 => "0000101011110010",
563 => "0000101011110100",564 => "0000101011110110",
565 => "0000101011110111",566 => "0000101011111001",
567 => "0000101011111011",568 => "0000101011111101",
569 => "0000101011111110",570 => "0000101100000000",
571 => "0000100001001101",572 => "0000101100000100",
573 => "0000101100000110",574 => "0000101100000111",
575 => "0000101100001001",576 => "0000101100001011",
577 => "0000101100001101",578 => "0000101100001110",
579 => "0000101100010000",580 => "0000101100010010",
581 => "0000101100010100",582 => "0000100001001111",
583 => "0000101100010111",584 => "0000101100011001",
585 => "0000101100011011",586 => "0000101100011101",
587 => "0000101100011111",588 => "0000100000001000",
589 => "0000101100100010",590 => "0000101100100100",
591 => "0000101100100110",592 => "0000101100101000",
593 => "0000101100101001",594 => "0000101100101011",
595 => "0000101100101101",596 => "0000101100101111",
597 => "0000101100110001",598 => "0000101100110010",
599 => "0000100001010010",600 => "0000101100110110",
601 => "0000101100111000",602 => "0000101100111010",
603 => "0000101100111100",604 => "0000101100111101",
605 => "0000101100111111",606 => "0000101101000001",
607 => "0000101101000011",608 => "0000101101000101",
609 => "0000101101000111",610 => "0000100001010100",
611 => "0000101101001010",612 => "0000101101001100",
613 => "0000101101001110",614 => "0000101101010000",
615 => "0000100001010101",616 => "0000101101010100",
617 => "0000101101010101",618 => "0000101101010111",
619 => "0000101101011001",620 => "0000101101011011",
621 => "0000101101011101",622 => "0000101101011111",
623 => "0000101101100001",624 => "0000101101100010",
625 => "0000101101100100",626 => "0000100001010111",
627 => "0000101101101000",628 => "0000101101101010",
629 => "0000101101101100",630 => "0000101101101110",
631 => "0000101101101111",632 => "0000101101110001",
633 => "0000101101110011",634 => "0000101101110101",
635 => "0000101101110111",636 => "0000101101111001",
637 => "0000101101111011",638 => "0000101101111101",
639 => "0000101101111111",640 => "0000101110000000",
641 => "0000101110000010",642 => "0000100000001001",
643 => "0000101110000110",644 => "0000101110001000",
645 => "0000101110001010",646 => "0000101110001100",
647 => "0000100001011011",648 => "0000101110010000",
649 => "0000101110010010",650 => "0000101110010100",
651 => "0000101110010101",652 => "0000101110010111",
653 => "0000101110011001",654 => "0000101110011011",
655 => "0000101110011101",656 => "0000101110011111",
657 => "0000101110100001",658 => "0000101110100011",
659 => "0000101110100101",660 => "0000101110100111",
661 => "0000101110101001",662 => "0000101110101011",
663 => "0000101110101101",664 => "0000101110101111",
665 => "0000101110110000",666 => "0000101110110010",
667 => "0000101110110100",668 => "0000100001011111",
669 => "0000101110111000",670 => "0000101110111010",
671 => "0000101110111100",672 => "0000101110111110",
673 => "0000100001100000",674 => "0000101111000010",
675 => "0000101111000100",676 => "0000101111000110",
677 => "0000101111001000",678 => "0000100001100001",
679 => "0000101111001100",680 => "0000101111001110",
681 => "0000101111010000",682 => "0000101111010010",
683 => "0000100001100010",684 => "0000101111010110",
685 => "0000101111011000",686 => "0000101111011010",
687 => "0000101111011100",688 => "0000100001100011",
689 => "0000101111100000",690 => "0000101111100010",
691 => "0000101111100100",692 => "0000101111100110",
693 => "0001000000000000",694 => "0001000000000010",
695 => "0001000000000100",696 => "0001000000000110",
697 => "0001000000001000",698 => "0001000000000001",
699 => "0001000000001100",700 => "0001000000001110",
701 => "0001000000010000",702 => "0001000000010010",
703 => "0001000000000010",704 => "0001000000010110",
705 => "0001000000011000",706 => "0001000000011010",
707 => "0001000000011100",708 => "0001000000000011",
709 => "0001000000100000",710 => "0001000000100010",
711 => "0001000000100100",712 => "0001000000100110",
713 => "0001000000000100",714 => "0001000000101010",
715 => "0001000000101100",716 => "0001000000101110",
717 => "0001000000110000",718 => "0001000000000101",
719 => "0001000000110100",720 => "0001000000110110",
721 => "0001000000111000",722 => "0001000000111011",
723 => "0001000000111101",724 => "0001000000111111",
725 => "0001000001000001",726 => "0001000001000011",
727 => "0001000001000101",728 => "0001000001000111",
729 => "0001000001001001",730 => "0001000001001011",
731 => "0001000001001101",732 => "0001000001001111",
733 => "0001000001010001",734 => "0001000001010011",
735 => "0001000001010101",736 => "0001000001011000",
737 => "0001000000001001",738 => "0001000001011100",
739 => "0001000001011110",740 => "0001000001100000",
741 => "0001000001100010",742 => "0001000000000001",
743 => "0001000001100110",744 => "0001000001101000",
745 => "0001000001101010",746 => "0001000001101101",
747 => "0001000001101111",748 => "0001000001110001",
749 => "0001000001110011",750 => "0001000001110101",
751 => "0001000001110111",752 => "0001000001111001",
753 => "0001000001111011",754 => "0001000001111101",
755 => "0001000010000000",756 => "0001000000001101",
757 => "0001000010000100",758 => "0001000010000110",
759 => "0001000010001000",760 => "0001000010001010",
761 => "0001000000001110",762 => "0001000010001111",
763 => "0001000010010001",764 => "0001000010010011",
765 => "0001000010010101",766 => "0001000010010111",
767 => "0001000010011001",768 => "0001000010011011",
769 => "0001000010011110",770 => "0001000000010000",
771 => "0001000010100010",772 => "0001000010100100",
773 => "0001000010100110",774 => "0001000010101000",
775 => "0001000010101011",776 => "0001000010101101",
777 => "0001000010101111",778 => "0001000010110001",
779 => "0001000010110011",780 => "0001000010110101",
781 => "0001000010111000",782 => "0001000010111010",
783 => "0001000010111100",784 => "0001000000010011",
785 => "0001000011000000",786 => "0001000011000011",
787 => "0001000011000101",788 => "0001000011000111",
789 => "0001000011001001",790 => "0001000011001011",
791 => "0001000011001110",792 => "0001000011010000",
793 => "0001000000010101",794 => "0001000011010100",
795 => "0001000011010110",796 => "0001000011011001",
797 => "0001000011011011",798 => "0001000011011101",
799 => "0001000011011111",800 => "0001000011100010",
801 => "0001000011100100",802 => "0001000000010111",
803 => "0001000011101000",804 => "0001000011101010",
805 => "0001000011101101",806 => "0001000011101111",
807 => "0001000011110001",808 => "0001000011110011",
809 => "0001000011110110",810 => "0001000011111000",
811 => "0001000000011001",812 => "0001000011111100",
813 => "0001000011111111",814 => "0001000100000001",
815 => "0001000100000011",816 => "0001000100000101",
817 => "0001000100001000",818 => "0001000100001010",
819 => "0001000100001100",820 => "0001000000011011",
821 => "0001000100010001",822 => "0001000100010011",
823 => "0001000100010101",824 => "0001000000011100",
825 => "0001000100011010",826 => "0001000100011100",
827 => "0001000100011110",828 => "0001000100100001",
829 => "0001000100100011",830 => "0001000100100101",
831 => "0001000100101000",832 => "0001000100101010",
833 => "0001000000000011",834 => "0001000100101111",
835 => "0001000100110001",836 => "0001000100110011",
837 => "0001000100110101",838 => "0001000100111000",
839 => "0001000100111010",840 => "0001000100111100",
841 => "0001000100111111",842 => "0001000101000001",
843 => "0001000101000011",844 => "0001000101000110",
845 => "0001000101001000",846 => "0001000000100001",
847 => "0001000101001101",848 => "0001000101001111",
849 => "0001000101010001",850 => "0001000000100010",
851 => "0001000101010110",852 => "0001000101011000",
853 => "0001000101011011",854 => "0001000101011101",
855 => "0001000101011111",856 => "0001000101100010",
857 => "0001000101100100",858 => "0001000101100110",
859 => "0001000101101001",860 => "0001000101101011",
861 => "0001000101101110",862 => "0001000101110000",
863 => "0001000000100101",864 => "0001000101110101",
865 => "0001000101110111",866 => "0001000101111001",
867 => "0001000000100110",868 => "0001000101111110",
869 => "0001000110000001",870 => "0001000110000011",
871 => "0001000110000101",872 => "0001000110001000",
873 => "0001000110001010",874 => "0001000110001100",
875 => "0001000110001111",876 => "0001000110010001",
877 => "0001000110010100",878 => "0001000110010110",
879 => "0001000110011000",880 => "0001000110011011",
881 => "0001000110011101",882 => "0001000110100000",
883 => "0001000110100010",884 => "0001000110100101",
885 => "0001000110100111",886 => "0001000110101001",
887 => "0001000110101100",888 => "0001000000101011",
889 => "0001000110110001",890 => "0001000110110011",
891 => "0001000110110110",892 => "0001000000101100",
893 => "0001000110111010",894 => "0001000110111101",
895 => "0001000110111111",896 => "0001000000101101",
897 => "0001000111000100",898 => "0001000111000111",
899 => "0001000111001001",900 => "0001000000101110",
901 => "0001000111001110",902 => "0001000111010001",
903 => "0001000111010011",904 => "0001000111010101",
905 => "0001000111011000",906 => "0001000111011010",
907 => "0001000111011101",908 => "0001000111011111",
909 => "0001000111100010",910 => "0001000111100100",
911 => "0001000111100111",912 => "0001000111101001",
913 => "0001000111101100",914 => "0001000111101110",
915 => "0001000111110001",916 => "0001000111110011",
917 => "0001000111110110",918 => "0001000111111000",
919 => "0001000111111011",920 => "0001000111111101",
921 => "0001001000000000",922 => "0001001000000010",
923 => "0001001000000101",924 => "0001001000000111",
925 => "0001001000001010",926 => "0001001000001100",
927 => "0001001000001111",928 => "0001001000010001",
929 => "0001001000010100",930 => "0001001000010111",
931 => "0001001000011001",932 => "0001000000110110",
933 => "0001001000011110",934 => "0001001000100001",
935 => "0001001000100011",936 => "0001000000110111",
937 => "0001001000101000",938 => "0001001000101011",
939 => "0001001000101101",940 => "0001000000111000",
941 => "0001001000110011",942 => "0001001000110101",
943 => "0001001000111000",944 => "0001000000111001",
945 => "0001001000111101",946 => "0001001000111111",
947 => "0001001001000010",948 => "0001001001000101",
949 => "0001001001000111",950 => "0001001001001010",
951 => "0001001001001100",952 => "0001001001001111",
953 => "0001001001010001",954 => "0001001001010100",
955 => "0001001001010111",956 => "0001001001011001",
957 => "0001001001011100",958 => "0001001001011110",
959 => "0001001001100001",960 => "0001001001100100",
961 => "0001001001100110",962 => "0001001001101001",
963 => "0001000000111110",964 => "0001001001101110",
965 => "0001001001110001",966 => "0001001001110011",
967 => "0001000000111111",968 => "0001001001111001",
969 => "0001001001111011",970 => "0001001001111110",
971 => "0001001010000001",972 => "0001001010000011",
973 => "0001001010000110",974 => "0001001010001001",
975 => "0001001010001011",976 => "0001001010001110",
977 => "0001001010010000",978 => "0001001010010011",
979 => "0001001010010110",980 => "0001001010011000",
981 => "0001001010011011",982 => "0001000001000011",
983 => "0001001010100000",984 => "0001001010100011",
985 => "0001001010100110",986 => "0001000001000100",
987 => "0001001010101011",988 => "0001001010101110",
989 => "0001001010110001",990 => "0001001010110011",
991 => "0001001010110110",992 => "0001001010111001",
993 => "0001001010111011",994 => "0001001010111110",
995 => "0001001011000001",996 => "0001001011000011",
997 => "0001000001000111",998 => "0001001011001001",
999 => "0001001011001100",1000 => "0000100001101001",
1001 => "0000100001101001",1002 => "0000100001101001",
1003 => "0000100001101010",1004 => "0000100001101010",
1005 => "0000100001101010",1006 => "0000100001101010",
1007 => "0000100001101010",1008 => "0000100001101010",
1009 => "0000100001101010",1010 => "0000100001101010",
1011 => "0000100001101010",1012 => "0000100001101010",
1013 => "0000100001101011",1014 => "0000100001101011",
1015 => "0000100001101011",1016 => "0000100001101011",
1017 => "0000100001101011",1018 => "0000100001101011",
1019 => "0000100001101011",1020 => "0000100001101011",
1021 => "0000100001101011",1022 => "0000100001101100",
1023 => "0000100001101100",1024 => "0000100001101100",
1025 => "0000100001101100",1026 => "0000100001101100",
1027 => "0000100001101100",1028 => "0000100001101100",
1029 => "0000100001101100",1030 => "0000100001101100",
1031 => "0000100001101101",1032 => "0000100001101101",
1033 => "0000100001101101",1034 => "0000100001101101",
1035 => "0000100001101101",1036 => "0000100001101101",
1037 => "0000100001101101",1038 => "0000100001101101",
1039 => "0000100001101101",1040 => "0000100000001011",
1041 => "0000100000001011",1042 => "0000100000001011",
1043 => "0000100000001011",1044 => "0000100000001011",
1045 => "0000100000001011",1046 => "0000100000001011",
1047 => "0000100000001011",1048 => "0000100000001011",
1049 => "0000100001101111",1050 => "0000100001101111",
1051 => "0000100001101111",1052 => "0000100001101111",
1053 => "0000100001101111",1054 => "0000100001101111",
1055 => "0000100001101111",1056 => "0000100001101111",
1057 => "0000100001101111",1058 => "0000100001110000",
1059 => "0000100001110000",1060 => "0000100001110000",
1061 => "0000100001110000",1062 => "0000100001110000",
1063 => "0000100001110000",1064 => "0000100001110000",
1065 => "0000100001110000",1066 => "0000100001110000",
1067 => "0000100001110001",1068 => "0000100001110001",
1069 => "0000100001110001",1070 => "0000100001110001",
1071 => "0000100001110001",1072 => "0000100001110001",
1073 => "0000100001110001",1074 => "0000100001110001",
1075 => "0000100001110001",1076 => "0000100001110010",
1077 => "0000100001110010",1078 => "0000100001110010",
1079 => "0000100001110010",1080 => "0000100001110010",
1081 => "0000100001110010",1082 => "0000100001110010",
1083 => "0000100001110010",1084 => "0000100001110010",
1085 => "0000100001110011",1086 => "0000100001110011",
1087 => "0000100001110011",1088 => "0000100001110011",
1089 => "0000100001110011",1090 => "0000100001110011",
1091 => "0000100001110011",1092 => "0000100001110011",
1093 => "0000100001110011",1094 => "0000100001110100",
1095 => "0000100001110100",1096 => "0000100001110100",
1097 => "0000100001110100",1098 => "0000100001110100",
1099 => "0000100001110100",1100 => "0000100001110100",
1101 => "0000100001110100",1102 => "0000100001110101",
1103 => "0000100001110101",1104 => "0000100001110101",
1105 => "0000100001110101",1106 => "0000100001110101",
1107 => "0000100001110101",1108 => "0000100001110101",
1109 => "0000100001110101",1110 => "0000100001110101",
1111 => "0000100001110110",1112 => "0000100001110110",
1113 => "0000100001110110",1114 => "0000100001110110",
1115 => "0000100001110110",1116 => "0000100001110110",
1117 => "0000100001110110",1118 => "0000100001110110",
1119 => "0000100001110110",1120 => "0000100001110111",
1121 => "0000100001110111",1122 => "0000100001110111",
1123 => "0000100001110111",1124 => "0000100001110111",
1125 => "0000100001110111",1126 => "0000100001110111",
1127 => "0000100001110111",1128 => "0000100001110111",
1129 => "0000100000001100",1130 => "0000100000001100",
1131 => "0000100000001100",1132 => "0000100000001100",
1133 => "0000100000001100",1134 => "0000100000001100",
1135 => "0000100000001100",1136 => "0000100000001100",
1137 => "0000100000001100",1138 => "0000100001111001",
1139 => "0000100001111001",1140 => "0000100001111001",
1141 => "0000100001111001",1142 => "0000100001111001",
1143 => "0000100001111001",1144 => "0000100001111001",
1145 => "0000100001111001",1146 => "0000100001111001",
1147 => "0000100001111010",1148 => "0000100001111010",
1149 => "0000100001111010",1150 => "0000100001111010",
1151 => "0000100001111010",1152 => "0000100001111010",
1153 => "0000100001111010",1154 => "0000100001111010",
1155 => "0000100001111010",1156 => "0000100001111011",
1157 => "0000100001111011",1158 => "0000100001111011",
1159 => "0000100001111011",1160 => "0000100001111011",
1161 => "0000100001111011",1162 => "0000100001111011",
1163 => "0000100001111011",1164 => "0000100001111011",
1165 => "0000100001111100",1166 => "0000100001111100",
1167 => "0000100001111100",1168 => "0000100001111100",
1169 => "0000100001111100",1170 => "0000100001111100",
1171 => "0000100001111100",1172 => "0000100001111100",
1173 => "0000100001111100",1174 => "0000100001111101",
1175 => "0000100001111101",1176 => "0000100001111101",
1177 => "0000100001111101",1178 => "0000100001111101",
1179 => "0000100001111101",1180 => "0000100001111101",
1181 => "0000100001111101",1182 => "0000100001111101",
1183 => "0000100001111110",1184 => "0000100001111110",
1185 => "0000100001111110",1186 => "0000100001111110",
1187 => "0000100001111110",1188 => "0000100001111110",
1189 => "0000100001111110",1190 => "0000100001111110",
1191 => "0000100001111110",1192 => "0000100001111111",
1193 => "0000100001111111",1194 => "0000100001111111",
1195 => "0000100001111111",1196 => "0000100001111111",
1197 => "0000100001111111",1198 => "0000100001111111",
1199 => "0000100001111111",1200 => "0000100001111111",
1201 => "0000100010000000",1202 => "0000100010000000",
1203 => "0000100010000000",1204 => "0000100010000000",
1205 => "0000100010000000",1206 => "0000100010000000",
1207 => "0000100010000000",1208 => "0000100010000000",
1209 => "0000100010000001",1210 => "0000100010000001",
1211 => "0000100010000001",1212 => "0000100010000001",
1213 => "0000100010000001",1214 => "0000100010000001",
1215 => "0000100010000001",1216 => "0000100010000001",
1217 => "0000100010000001",1218 => "0000100000001101",
1219 => "0000100000001101",1220 => "0000100000001101",
1221 => "0000100000001101",1222 => "0000100000001101",
1223 => "0000100000001101",1224 => "0000100000001101",
1225 => "0000100000001101",1226 => "0000100000001101",
1227 => "0000100010000011",1228 => "0000100010000011",
1229 => "0000100010000011",1230 => "0000100010000011",
1231 => "0000100010000011",1232 => "0000100010000011",
1233 => "0000100010000011",1234 => "0000100010000011",
1235 => "0000100010000011",1236 => "0000100010000100",
1237 => "0000100010000100",1238 => "0000100010000100",
1239 => "0000100010000100",1240 => "0000100010000100",
1241 => "0000100010000100",1242 => "0000100010000100",
1243 => "0000100010000100",1244 => "0000100010000100",
1245 => "0000100010000101",1246 => "0000100010000101",
1247 => "0000100010000101",1248 => "0000100010000101",
1249 => "0000100010000101",1250 => "0000100010000101",
1251 => "0000100010000101",1252 => "0000100010000101",
1253 => "0000100010000101",1254 => "0000100010000110",
1255 => "0000100010000110",1256 => "0000100010000110",
1257 => "0000100010000110",1258 => "0000100010000110",
1259 => "0000100010000110",1260 => "0000100010000110",
1261 => "0000100010000110",1262 => "0000100010000111",
1263 => "0000100010000111",1264 => "0000100010000111",
1265 => "0000100010000111",1266 => "0000100010000111",
1267 => "0000100010000111",1268 => "0000100010000111",
1269 => "0000100010000111",1270 => "0000100010000111",
1271 => "0000100010001000",1272 => "0000100010001000",
1273 => "0000100010001000",1274 => "0000100010001000",
1275 => "0000100010001000",1276 => "0000100010001000",
1277 => "0000100010001000",1278 => "0000100010001000",
1279 => "0000100010001000",1280 => "0000100010001001",
1281 => "0000100010001001",1282 => "0000100010001001",
1283 => "0000100010001001",1284 => "0000100010001001",
1285 => "0000100010001001",1286 => "0000100010001001",
1287 => "0000100010001001",1288 => "0000100010001001",
1289 => "0000100010001010",1290 => "0000100010001010",
1291 => "0000100010001010",1292 => "0000100010001010",
1293 => "0000100010001010",1294 => "0000100010001010",
1295 => "0000100010001010",1296 => "0000100010001010",
1297 => "0000100010001010",1298 => "0000100010001011",
1299 => "0000100010001011",1300 => "0000100010001011",
1301 => "0000100010001011",1302 => "0000100010001011",
1303 => "0000100010001011",1304 => "0000100010001011",
1305 => "0000100010001011",1306 => "0000100000001110",
1307 => "0000100000001110",1308 => "0000100000001110",
1309 => "0000100000001110",1310 => "0000100000001110",
1311 => "0000100000001110",1312 => "0000100000001110",
1313 => "0000100000001110",1314 => "0000100000001110",
1315 => "0000100010001101",1316 => "0000100010001101",
1317 => "0000100010001101",1318 => "0000100010001101",
1319 => "0000100010001101",1320 => "0000100010001101",
1321 => "0000100010001101",1322 => "0000100010001101",
1323 => "0000100010001101",1324 => "0000100010001110",
1325 => "0000100010001110",1326 => "0000100010001110",
1327 => "0000100010001110",1328 => "0000100010001110",
1329 => "0000100010001110",1330 => "0000100010001110",
1331 => "0000100010001110",1332 => "0000100010001110",
1333 => "0000100010001111",1334 => "0000100010001111",
1335 => "0000100010001111",1336 => "0000100010001111",
1337 => "0000100010001111",1338 => "0000100010001111",
1339 => "0000100010001111",1340 => "0000100010001111",
1341 => "0000100010010000",1342 => "0000100010010000",
1343 => "0000100010010000",1344 => "0000100010010000",
1345 => "0000100010010000",1346 => "0000100010010000",
1347 => "0000100010010000",1348 => "0000100010010000",
1349 => "0000100010010000",1350 => "0000100010010001",
1351 => "0000100010010001",1352 => "0000100010010001",
1353 => "0000100010010001",1354 => "0000100010010001",
1355 => "0000100010010001",1356 => "0000100010010001",
1357 => "0000100010010001",1358 => "0000100010010001",
1359 => "0000100010010010",1360 => "0000100010010010",
1361 => "0000100010010010",1362 => "0000100010010010",
1363 => "0000100010010010",1364 => "0000100010010010",
1365 => "0000100010010010",1366 => "0000100010010010",
1367 => "0000100010010010",1368 => "0000100010010011",
1369 => "0000100010010011",1370 => "0000100010010011",
1371 => "0000100010010011",1372 => "0000100010010011",
1373 => "0000100010010011",1374 => "0000100010010011",
1375 => "0000100010010011",1376 => "0000100010010100",
1377 => "0000100010010100",1378 => "0000100010010100",
1379 => "0000100010010100",1380 => "0000100010010100",
1381 => "0000100010010100",1382 => "0000100010010100",
1383 => "0000100010010100",1384 => "0000100010010100",
1385 => "0000100010010101",1386 => "0000100010010101",
1387 => "0000100010010101",1388 => "0000100010010101",
1389 => "0000100010010101",1390 => "0000100010010101",
1391 => "0000100010010101",1392 => "0000100010010101",
1393 => "0000100010010101",1394 => "0000100000001111",
1395 => "0000100000001111",1396 => "0000100000001111",
1397 => "0000100000001111",1398 => "0000100000001111",
1399 => "0000100000001111",1400 => "0000100000001111",
1401 => "0000100000001111",1402 => "0000100010010111",
1403 => "0000100010010111",1404 => "0000100010010111",
1405 => "0000100010010111",1406 => "0000100010010111",
1407 => "0000100010010111",1408 => "0000100010010111",
1409 => "0000100010010111",1410 => "0000100010010111",
1411 => "0000100010011000",1412 => "0000100010011000",
1413 => "0000100010011000",1414 => "0000100010011000",
1415 => "0000100010011000",1416 => "0000100010011000",
1417 => "0000100010011000",1418 => "0000100010011000",
1419 => "0000100010011000",1420 => "0000100010011001",
1421 => "0000100010011001",1422 => "0000100010011001",
1423 => "0000100010011001",1424 => "0000100010011001",
1425 => "0000100010011001",1426 => "0000100010011001",
1427 => "0000100010011001",1428 => "0000100010011001",
1429 => "0000100010011010",1430 => "0000100010011010",
1431 => "0000100010011010",1432 => "0000100010011010",
1433 => "0000100010011010",1434 => "0000100010011010",
1435 => "0000100010011010",1436 => "0000100010011010",
1437 => "0000100010011011",1438 => "0000100010011011",
1439 => "0000100010011011",1440 => "0000100010011011",
1441 => "0000100010011011",1442 => "0000100010011011",
1443 => "0000100010011011",1444 => "0000100010011011",
1445 => "0000100010011011",1446 => "0000100010011100",
1447 => "0000100010011100",1448 => "0000100010011100",
1449 => "0000100010011100",1450 => "0000100010011100",
1451 => "0000100010011100",1452 => "0000100010011100",
1453 => "0000100010011100",1454 => "0000100010011101",
1455 => "0000100010011101",1456 => "0000100010011101",
1457 => "0000100010011101",1458 => "0000100010011101",
1459 => "0000100010011101",1460 => "0000100010011101",
1461 => "0000100010011101",1462 => "0000100010011101",
1463 => "0000100010011110",1464 => "0000100010011110",
1465 => "0000100010011110",1466 => "0000100010011110",
1467 => "0000100010011110",1468 => "0000100010011110",
1469 => "0000100010011110",1470 => "0000100010011110",
1471 => "0000100010011110",1472 => "0000100010011111",
1473 => "0000100010011111",1474 => "0000100010011111",
1475 => "0000100010011111",1476 => "0000100010011111",
1477 => "0000100010011111",1478 => "0000100010011111",
1479 => "0000100010011111",1480 => "0000100000010000",
1481 => "0000100000010000",1482 => "0000100000010000",
1483 => "0000100000010000",1484 => "0000100000010000",
1485 => "0000100000010000",1486 => "0000100000010000",
1487 => "0000100000010000",1488 => "0000100000010000",
1489 => "0000100010100001",1490 => "0000100010100001",
1491 => "0000100010100001",1492 => "0000100010100001",
1493 => "0000100010100001",1494 => "0000100010100001",
1495 => "0000100010100001",1496 => "0000100010100001",
1497 => "0000100010100001",1498 => "0000100010100010",
1499 => "0000100010100010",1500 => "0000100010100010",
1501 => "0000100010100010",1502 => "0000100010100010",
1503 => "0000100010100010",1504 => "0000100010100010",
1505 => "0000100010100010",1506 => "0000100010100011",
1507 => "0000100010100011",1508 => "0000100010100011",
1509 => "0000100010100011",1510 => "0000100010100011",
1511 => "0000100010100011",1512 => "0000100010100011",
1513 => "0000100010100011",1514 => "0000100010100011",
1515 => "0000100010100100",1516 => "0000100010100100",
1517 => "0000100010100100",1518 => "0000100010100100",
1519 => "0000100010100100",1520 => "0000100010100100",
1521 => "0000100010100100",1522 => "0000100010100100",
1523 => "0000100010100101",1524 => "0000100010100101",
1525 => "0000100010100101",1526 => "0000100010100101",
1527 => "0000100010100101",1528 => "0000100010100101",
1529 => "0000100010100101",1530 => "0000100010100101",
1531 => "0000100010100101",1532 => "0000100010100110",
1533 => "0000100010100110",1534 => "0000100010100110",
1535 => "0000100010100110",1536 => "0000100010100110",
1537 => "0000100010100110",1538 => "0000100010100110",
1539 => "0000100010100110",1540 => "0000100010100110",
1541 => "0000100010100111",1542 => "0000100010100111",
1543 => "0000100010100111",1544 => "0000100010100111",
1545 => "0000100010100111",1546 => "0000100010100111",
1547 => "0000100010100111",1548 => "0000100010100111",
1549 => "0000100010101000",1550 => "0000100010101000",
1551 => "0000100010101000",1552 => "0000100010101000",
1553 => "0000100010101000",1554 => "0000100010101000",
1555 => "0000100010101000",1556 => "0000100010101000",
1557 => "0000100010101000",1558 => "0000100010101001",
1559 => "0000100010101001",1560 => "0000100010101001",
1561 => "0000100010101001",1562 => "0000100010101001",
1563 => "0000100010101001",1564 => "0000100010101001",
1565 => "0000100010101001",1566 => "0000100000010001",
1567 => "0000100000010001",1568 => "0000100000010001",
1569 => "0000100000010001",1570 => "0000100000010001",
1571 => "0000100000010001",1572 => "0000100000010001",
1573 => "0000100000010001",1574 => "0000100000010001",
1575 => "0000100010101011",1576 => "0000100010101011",
1577 => "0000100010101011",1578 => "0000100010101011",
1579 => "0000100010101011",1580 => "0000100010101011",
1581 => "0000100010101011",1582 => "0000100010101011",
1583 => "0000100010101100",1584 => "0000100010101100",
1585 => "0000100010101100",1586 => "0000100010101100",
1587 => "0000100010101100",1588 => "0000100010101100",
1589 => "0000100010101100",1590 => "0000100010101100",
1591 => "0000100010101100",1592 => "0000100010101101",
1593 => "0000100010101101",1594 => "0000100010101101",
1595 => "0000100010101101",1596 => "0000100010101101",
1597 => "0000100010101101",1598 => "0000100010101101",
1599 => "0000100010101101",1600 => "0000100010101110",
1601 => "0000100010101110",1602 => "0000100010101110",
1603 => "0000100010101110",1604 => "0000100010101110",
1605 => "0000100010101110",1606 => "0000100010101110",
1607 => "0000100010101110",1608 => "0000100010101110",
1609 => "0000100010101111",1610 => "0000100010101111",
1611 => "0000100010101111",1612 => "0000100010101111",
1613 => "0000100010101111",1614 => "0000100010101111",
1615 => "0000100010101111",1616 => "0000100010101111",
1617 => "0000100010110000",1618 => "0000100010110000",
1619 => "0000100010110000",1620 => "0000100010110000",
1621 => "0000100010110000",1622 => "0000100010110000",
1623 => "0000100010110000",1624 => "0000100010110000",
1625 => "0000100010110000",1626 => "0000100010110001",
1627 => "0000100010110001",1628 => "0000100010110001",
1629 => "0000100010110001",1630 => "0000100010110001",
1631 => "0000100010110001",1632 => "0000100010110001",
1633 => "0000100010110001",1634 => "0000100010110010",
1635 => "0000100010110010",1636 => "0000100010110010",
1637 => "0000100010110010",1638 => "0000100010110010",
1639 => "0000100010110010",1640 => "0000100010110010",
1641 => "0000100010110010",1642 => "0000100010110010",
1643 => "0000100010110011",1644 => "0000100010110011",
1645 => "0000100010110011",1646 => "0000100010110011",
1647 => "0000100010110011",1648 => "0000100010110011",
1649 => "0000100010110011",1650 => "0000100010110011",
1651 => "0000100000010010",1652 => "0000100000010010",
1653 => "0000100000010010",1654 => "0000100000010010",
1655 => "0000100000010010",1656 => "0000100000010010",
1657 => "0000100000010010",1658 => "0000100000010010",
1659 => "0000100000010010",1660 => "0000100010110101",
1661 => "0000100010110101",1662 => "0000100010110101",
1663 => "0000100010110101",1664 => "0000100010110101",
1665 => "0000100010110101",1666 => "0000100010110101",
1667 => "0000100010110101",1668 => "0000100010110110",
1669 => "0000100010110110",1670 => "0000100010110110",
1671 => "0000100010110110",1672 => "0000100010110110",
1673 => "0000100010110110",1674 => "0000100010110110",
1675 => "0000100010110110",1676 => "0000100010110110",
1677 => "0000100010110111",1678 => "0000100010110111",
1679 => "0000100010110111",1680 => "0000100010110111",
1681 => "0000100010110111",1682 => "0000100010110111",
1683 => "0000100010110111",1684 => "0000100010110111",
1685 => "0000100010111000",1686 => "0000100010111000",
1687 => "0000100010111000",1688 => "0000100010111000",
1689 => "0000100010111000",1690 => "0000100010111000",
1691 => "0000100010111000",1692 => "0000100010111000",
1693 => "0000100010111000",1694 => "0000100010111001",
1695 => "0000100010111001",1696 => "0000100010111001",
1697 => "0000100010111001",1698 => "0000100010111001",
1699 => "0000100010111001",1700 => "0000100010111001",
1701 => "0000100010111001",1702 => "0000100010111010",
1703 => "0000100010111010",1704 => "0000100010111010",
1705 => "0000100010111010",1706 => "0000100010111010",
1707 => "0000100010111010",1708 => "0000100010111010",
1709 => "0000100010111010",1710 => "0000100010111010",
1711 => "0000100010111011",1712 => "0000100010111011",
1713 => "0000100010111011",1714 => "0000100010111011",
1715 => "0000100010111011",1716 => "0000100010111011",
1717 => "0000100010111011",1718 => "0000100010111011",
1719 => "0000100010111100",1720 => "0000100010111100",
1721 => "0000100010111100",1722 => "0000100010111100",
1723 => "0000100010111100",1724 => "0000100010111100",
1725 => "0000100010111100",1726 => "0000100010111100",
1727 => "0000100010111101",1728 => "0000100010111101",
1729 => "0000100010111101",1730 => "0000100010111101",
1731 => "0000100010111101",1732 => "0000100010111101",
1733 => "0000100010111101",1734 => "0000100010111101",
1735 => "0000100010111101",1736 => "0000100000010011",
1737 => "0000100000010011",1738 => "0000100000010011",
1739 => "0000100000010011",1740 => "0000100000010011",
1741 => "0000100000010011",1742 => "0000100000010011",
1743 => "0000100000010011",1744 => "0000100010111111",
1745 => "0000100010111111",1746 => "0000100010111111",
1747 => "0000100010111111",1748 => "0000100010111111",
1749 => "0000100010111111",1750 => "0000100010111111",
1751 => "0000100010111111",1752 => "0000100010111111",
1753 => "0000100011000000",1754 => "0000100011000000",
1755 => "0000100011000000",1756 => "0000100011000000",
1757 => "0000100011000000",1758 => "0000100011000000",
1759 => "0000100011000000",1760 => "0000100011000000",
1761 => "0000100011000001",1762 => "0000100011000001",
1763 => "0000100011000001",1764 => "0000100011000001",
1765 => "0000100011000001",1766 => "0000100011000001",
1767 => "0000100011000001",1768 => "0000100011000001",
1769 => "0000100011000010",1770 => "0000100011000010",
1771 => "0000100011000010",1772 => "0000100011000010",
1773 => "0000100011000010",1774 => "0000100011000010",
1775 => "0000100011000010",1776 => "0000100011000010",
1777 => "0000100011000010",1778 => "0000100011000011",
1779 => "0000100011000011",1780 => "0000100011000011",
1781 => "0000100011000011",1782 => "0000100011000011",
1783 => "0000100011000011",1784 => "0000100011000011",
1785 => "0000100011000011",1786 => "0000100011000100",
1787 => "0000100011000100",1788 => "0000100011000100",
1789 => "0000100011000100",1790 => "0000100011000100",
1791 => "0000100011000100",1792 => "0000100011000100",
1793 => "0000100011000100",1794 => "0000100011000100",
1795 => "0000100011000101",1796 => "0000100011000101",
1797 => "0000100011000101",1798 => "0000100011000101",
1799 => "0000100011000101",1800 => "0000100011000101",
1801 => "0000100011000101",1802 => "0000100011000101",
1803 => "0000100011000110",1804 => "0000100011000110",
1805 => "0000100011000110",1806 => "0000100011000110",
1807 => "0000100011000110",1808 => "0000100011000110",
1809 => "0000100011000110",1810 => "0000100011000110",
1811 => "0000100011000111",1812 => "0000100011000111",
1813 => "0000100011000111",1814 => "0000100011000111",
1815 => "0000100011000111",1816 => "0000100011000111",
1817 => "0000100011000111",1818 => "0000100011000111",
1819 => "0000100011000111",1820 => "0000100000000010",
1821 => "0000100000000010",1822 => "0000100000000010",
1823 => "0000100000000010",1824 => "0000100000000010",
1825 => "0000100000000010",1826 => "0000100000000010",
1827 => "0000100000000010",1828 => "0000100011001001",
1829 => "0000100011001001",1830 => "0000100011001001",
1831 => "0000100011001001",1832 => "0000100011001001",
1833 => "0000100011001001",1834 => "0000100011001001",
1835 => "0000100011001001",1836 => "0000100011001010",
1837 => "0000100011001010",1838 => "0000100011001010",
1839 => "0000100011001010",1840 => "0000100011001010",
1841 => "0000100011001010",1842 => "0000100011001010",
1843 => "0000100011001010",1844 => "0000100011001010",
1845 => "0000100011001011",1846 => "0000100011001011",
1847 => "0000100011001011",1848 => "0000100011001011",
1849 => "0000100011001011",1850 => "0000100011001011",
1851 => "0000100011001011",1852 => "0000100011001011",
1853 => "0000100011001100",1854 => "0000100011001100",
1855 => "0000100011001100",1856 => "0000100011001100",
1857 => "0000100011001100",1858 => "0000100011001100",
1859 => "0000100011001100",1860 => "0000100011001100",
1861 => "0000100011001101",1862 => "0000100011001101",
1863 => "0000100011001101",1864 => "0000100011001101",
1865 => "0000100011001101",1866 => "0000100011001101",
1867 => "0000100011001101",1868 => "0000100011001101",
1869 => "0000100011001110",1870 => "0000100011001110",
1871 => "0000100011001110",1872 => "0000100011001110",
1873 => "0000100011001110",1874 => "0000100011001110",
1875 => "0000100011001110",1876 => "0000100011001110",
1877 => "0000100011001110",1878 => "0000100011001111",
1879 => "0000100011001111",1880 => "0000100011001111",
1881 => "0000100011001111",1882 => "0000100011001111",
1883 => "0000100011001111",1884 => "0000100011001111",
1885 => "0000100011001111",1886 => "0000100011010000",
1887 => "0000100011010000",1888 => "0000100011010000",
1889 => "0000100011010000",1890 => "0000100011010000",
1891 => "0000100011010000",1892 => "0000100011010000",
1893 => "0000100011010000",1894 => "0000100011010001",
1895 => "0000100011010001",1896 => "0000100011010001",
1897 => "0000100011010001",1898 => "0000100011010001",
1899 => "0000100011010001",1900 => "0000100011010001",
1901 => "0000100011010001",1902 => "0000100011010001",
1903 => "0000100000010101",1904 => "0000100000010101",
1905 => "0000100000010101",1906 => "0000100000010101",
1907 => "0000100000010101",1908 => "0000100000010101",
1909 => "0000100000010101",1910 => "0000100000010101",
1911 => "0000100011010011",1912 => "0000100011010011",
1913 => "0000100011010011",1914 => "0000100011010011",
1915 => "0000100011010011",1916 => "0000100011010011",
1917 => "0000100011010011",1918 => "0000100011010011",
1919 => "0000100011010100",1920 => "0000100011010100",
1921 => "0000100011010100",1922 => "0000100011010100",
1923 => "0000100011010100",1924 => "0000100011010100",
1925 => "0000100011010100",1926 => "0000100011010100",
1927 => "0000100011010101",1928 => "0000100011010101",
1929 => "0000100011010101",1930 => "0000100011010101",
1931 => "0000100011010101",1932 => "0000100011010101",
1933 => "0000100011010101",1934 => "0000100011010101",
1935 => "0000100011010101",1936 => "0000100011010110",
1937 => "0000100011010110",1938 => "0000100011010110",
1939 => "0000100011010110",1940 => "0000100011010110",
1941 => "0000100011010110",1942 => "0000100011010110",
1943 => "0000100011010110",1944 => "0000100011010111",
1945 => "0000100011010111",1946 => "0000100011010111",
1947 => "0000100011010111",1948 => "0000100011010111",
1949 => "0000100011010111",1950 => "0000100011010111",
1951 => "0000100011010111",1952 => "0000100011011000",
1953 => "0000100011011000",1954 => "0000100011011000",
1955 => "0000100011011000",1956 => "0000100011011000",
1957 => "0000100011011000",1958 => "0000100011011000",
1959 => "0000100011011000",1960 => "0000100011011001",
1961 => "0000100011011001",1962 => "0000100011011001",
1963 => "0000100011011001",1964 => "0000100011011001",
1965 => "0000100011011001",1966 => "0000100011011001",
1967 => "0000100011011001",1968 => "0000100011011010",
1969 => "0000100011011010",1970 => "0000100011011010",
1971 => "0000100011011010",1972 => "0000100011011010",
1973 => "0000100011011010",1974 => "0000100011011010",
1975 => "0000100011011010",1976 => "0000100011011010",
1977 => "0000100011011011",1978 => "0000100011011011",
1979 => "0000100011011011",1980 => "0000100011011011",
1981 => "0000100011011011",1982 => "0000100011011011",
1983 => "0000100011011011",1984 => "0000100011011011",
1985 => "0000100000010110",1986 => "0000100000010110",
1987 => "0000100000010110",1988 => "0000100000010110",
1989 => "0000100000010110",1990 => "0000100000010110",
1991 => "0000100000010110",1992 => "0000100000010110",
1993 => "0000100011011101",1994 => "0000100011011101",
1995 => "0000100011011101",1996 => "0000100011011101",
1997 => "0000100011011101",1998 => "0000100011011101",
1999 => "0000100011011101",2000 => "0000100011011101",
2001 => "0000100011011110",2002 => "0000100011011110",
2003 => "0000100011011110",2004 => "0000100011011110",
2005 => "0000100011011110",2006 => "0000100011011110",
2007 => "0000100011011110",2008 => "0000100011011110",
2009 => "0000100011011111",2010 => "0000100011011111",
2011 => "0000100011011111",2012 => "0000100011011111",
2013 => "0000100011011111",2014 => "0000100011011111",
2015 => "0000100011011111",2016 => "0000100011011111",
2017 => "0000100011011111",2018 => "0000100011100000",
2019 => "0000100011100000",2020 => "0000100011100000",
2021 => "0000100011100000",2022 => "0000100011100000",
2023 => "0000100011100000",2024 => "0000100011100000",
2025 => "0000100011100000",2026 => "0000100011100001",
2027 => "0000100011100001",2028 => "0000100011100001",
2029 => "0000100011100001",2030 => "0000100011100001",
2031 => "0000100011100001",2032 => "0000100011100001",
2033 => "0000100011100001",2034 => "0000100011100010",
2035 => "0000100011100010",2036 => "0000100011100010",
2037 => "0000100011100010",2038 => "0000100011100010",
2039 => "0000100011100010",2040 => "0000100011100010",
2041 => "0000100011100010",2042 => "0000100011100011",
2043 => "0000100011100011",2044 => "0000100011100011",
2045 => "0000100011100011",2046 => "0000100011100011",
2047 => "0000100011100011",2048 => "0001001011001110",
2049 => "0001100000000100",2050 => "0001100000100000",
2051 => "0001101010011101",2052 => "0010000000110111",
2053 => "0010000111100010",2054 => "0010001110111001",
2055 => "0010100111011010",2056 => "0011000000000101",
2057 => "0011001010101110",2058 => "0001100000000100",
2059 => "0001100000100010",2060 => "0001100001000001",
2061 => "0001100001100000",2062 => "0001100001111111",
2063 => "0001100010011110",2064 => "0001100000010011",
2065 => "0001100011011110",2066 => "0001100011111110",
2067 => "0001100100011111",2068 => "0001100000100000",
2069 => "0001100101100001",2070 => "0001100110000011",
2071 => "0001100110100101",2072 => "0001100111001000",
2073 => "0001100000110001",2074 => "0001101000001101",
2075 => "0001101000110001",2076 => "0001101001010101",
2077 => "0001101001111001",2078 => "0001101010011101",
2079 => "0001101011000010",2080 => "0001101011100111",
2081 => "0001101100001101",2082 => "0001101100110011",
2083 => "0001101101011001",2084 => "0001101110000000",
2085 => "0001101110100111",2086 => "0001101111001111",
2087 => "0010000000001111",2088 => "0010000000110111",
2089 => "0010000001100000",2090 => "0010000010001001",
2091 => "0010000010110011",2092 => "0010000011011101",
2093 => "0010000100000111",2094 => "0010000100110010",
2095 => "0010000101011101",2096 => "0010000110001001",
2097 => "0010000110110101",2098 => "0010000111100010",
2099 => "0010001000001111",2100 => "0010001000111100",
2101 => "0010001001101010",2102 => "0010001010011001",
2103 => "0010001011000111",2104 => "0010001011110111",
2105 => "0010001100100111",2106 => "0010001101010111",
2107 => "0010001110001000",2108 => "0010001110111001",
2109 => "0010100000000011",2110 => "0010100000110101",
2111 => "0010100001101000",2112 => "0010100010011011",
2113 => "0010100011001111",2114 => "0010100100000011",
2115 => "0010100100111000",2116 => "0010100101101110",
2117 => "0010100110100011",2118 => "0010100111011010",
2119 => "0010101000010001",2120 => "0010101001001001",
2121 => "0010101010000001",2122 => "0010101010111001",
2123 => "0010101011110011",2124 => "0010101100101100",
2125 => "0010101101100111",2126 => "0010100001011101",
2127 => "0010101111011101",2128 => "0011000000000101",
2129 => "0011000000001011",2130 => "0011000010101100",
2131 => "0011000011101010",2132 => "0011000100101001",
2133 => "0011000000100100",2134 => "0011000110101000",
2135 => "0011000111101000",2136 => "0011001000101010",
2137 => "0011001001101011",2138 => "0011001010101110",
2139 => "0011001011110001",2140 => "0011001100110101",
2141 => "0011000001011001",2142 => "0011001110111111",
2143 => "0011100000011101",2144 => "0011100001100011",
2145 => "0011100010101011",2146 => "0011100011110011",
2147 => "0011100100111100",2148 => "0001100000000100",
2149 => "0001100000000111",2150 => "0001100000000001",
2151 => "0001100000001101",2152 => "0001100000010000",
2153 => "0001100000010011",2154 => "0001100000010110",
2155 => "0001100000011001",2156 => "0001100000011100",
2157 => "0001100000011111",2158 => "0001100000100010",
2159 => "0001100000100101",2160 => "0001100000000100",
2161 => "0001100000101011",2162 => "0001100000101111",
2163 => "0001100000000101",2164 => "0001100000110101",
2165 => "0001100000111000",2166 => "0001100000111011",
2167 => "0001100000111110",2168 => "0001100001000001",
2169 => "0001100001000100",2170 => "0001100001000111",
2171 => "0001100001001010",2172 => "0001100001001101",
2173 => "0001100000001000",2174 => "0001100001010011",
2175 => "0001100001010110",2176 => "0001100001011001",
2177 => "0001100001011101",2178 => "0001100001100000",
2179 => "0001100001100011",2180 => "0001100001100110",
2181 => "0001100001101001",2182 => "0001100001101100",
2183 => "0001100001101111",2184 => "0001100001110010",
2185 => "0001100001110101",2186 => "0001100001111001",
2187 => "0001100001111100",2188 => "0001100001111111",
2189 => "0001100000001101",2190 => "0001100010000101",
2191 => "0001100010001000",2192 => "0001100010001011",
2193 => "0001100010001110",2194 => "0001100010010010",
2195 => "0001100010010101",2196 => "0001100010011000",
2197 => "0001100010011011",2198 => "0001100010011110",
2199 => "0001100010100001",2200 => "0001100010100101",
2201 => "0001100010101000",2202 => "0001100010101011",
2203 => "0001100010101110",2204 => "0001100010110001",
2205 => "0001100000010010",2206 => "0001100010111000",
2207 => "0001100010111011",2208 => "0001100000010011",
2209 => "0001100011000001",2210 => "0001100011000100",
2211 => "0001100000000010",2212 => "0001100011001011",
2213 => "0001100011001110",2214 => "0001100011010001",
2215 => "0001100011010100",2216 => "0001100011011000",
2217 => "0001100011011011",2218 => "0001100011011110",
2219 => "0001100011100001",2220 => "0001100011100100",
2221 => "0001100011101000",2222 => "0001100011101011",
2223 => "0001100011101110",2224 => "0001100011110001",
2225 => "0001100011110101",2226 => "0001100011111000",
2227 => "0001100011111011",2228 => "0001100011111110",
2229 => "0001100100000010",2230 => "0001100100000101",
2231 => "0001100100001000",2232 => "0001100100001011",
2233 => "0001100100001111",2234 => "0001100100010010",
2235 => "0001100100010101",2236 => "0001100100011001",
2237 => "0001100100011100",2238 => "0001100100011111",
2239 => "0001100000011101",2240 => "0001100100100110",
2241 => "0001100100101001",2242 => "0001100000000011",
2243 => "0001100100110000",2244 => "0001100100110011",
2245 => "0001100000011111",2246 => "0001100100111001",
2247 => "0001100100111101",2248 => "0001100000100000",
2249 => "0001100101000011",2250 => "0001100101000111",
2251 => "0001100000100001",2252 => "0001100101001101",
2253 => "0001100101010001",2254 => "0001100000100010",
2255 => "0001100101010111",2256 => "0001100101011011",
2257 => "0001100000100011",2258 => "0001100101100001",
2259 => "0001100101100101",2260 => "0001100000100100",
2261 => "0001100101101100",2262 => "0001100101101111",
2263 => "0001100000100101",2264 => "0001100101110110",
2265 => "0001100101111001",2266 => "0001100000100110",
2267 => "0001100110000000",2268 => "0001100110000011",
2269 => "0001100110000111",2270 => "0001100110001010",
2271 => "0001100110001101",2272 => "0001100110010001",
2273 => "0001100110010100",2274 => "0001100110011000",
2275 => "0001100110011011",2276 => "0001100110011110",
2277 => "0001100110100010",2278 => "0001100110100101",
2279 => "0001100110101001",2280 => "0001100110101100",
2281 => "0001100110110000",2282 => "0001100110110011",
2283 => "0001100110110110",2284 => "0001100110111010",
2285 => "0001100110111101",2286 => "0001100111000001",
2287 => "0001100111000100",2288 => "0001100111001000",
2289 => "0001100111001011",2290 => "0001100111001111",
2291 => "0001100111010010",2292 => "0001100111010101",
2293 => "0001100111011001",2294 => "0001100111011100",
2295 => "0001100000110000",2296 => "0001100111100011",
2297 => "0001100111100111",2298 => "0001100000110001",
2299 => "0001100111101110",2300 => "0001100111110001",
2301 => "0001100111110101",2302 => "0001100111111000",
2303 => "0001100111111100",2304 => "0001100111111111",
2305 => "0001101000000011",2306 => "0001101000000110",
2307 => "0001101000001010",2308 => "0001101000001101",
2309 => "0001101000010001",2310 => "0001101000010100",
2311 => "0001101000011000",2312 => "0001100000110110",
2313 => "0001101000011111",2314 => "0001101000100011",
2315 => "0001100000110111",2316 => "0001101000101010",
2317 => "0001101000101101",2318 => "0001101000110001",
2319 => "0001101000110100",2320 => "0001101000111000",
2321 => "0001101000111100",2322 => "0001101000111111",
2323 => "0001101001000011",2324 => "0001101001000110",
2325 => "0001101001001010",2326 => "0001101001001101",
2327 => "0001101001010001",2328 => "0001101001010101",
2329 => "0001100000000110",2330 => "0001101001011100",
2331 => "0001101001011111",2332 => "0001101001100011",
2333 => "0001101001100111",2334 => "0001101001101010",
2335 => "0001101001101110",2336 => "0001101001110010",
2337 => "0001101001110101",2338 => "0001101001111001",
2339 => "0001101001111100",2340 => "0001100001000000",
2341 => "0001101010000100",2342 => "0001101010000111",
2343 => "0001101010001011",2344 => "0001101010001111",
2345 => "0001101010010010",2346 => "0001101010010110",
2347 => "0001101010011010",2348 => "0001101010011101",
2349 => "0001101010100001",2350 => "0001101010100101",
2351 => "0001100001000100",2352 => "0001101010101100",
2353 => "0001101010110000",2354 => "0001101010110011",
2355 => "0001101010110111",2356 => "0001101010111011",
2357 => "0001101010111110",2358 => "0001101011000010",
2359 => "0001100001000111",2360 => "0001101011001010",
2361 => "0001101011001101",2362 => "0001101011010001",
2363 => "0001101011010101",2364 => "0001101011011000",
2365 => "0001101011011100",2366 => "0001101011100000",
2367 => "0001100001001010",2368 => "0001101011100111",
2369 => "0001101011101011",2370 => "0001101011101111",
2371 => "0001101011110011",2372 => "0001101011110110",
2373 => "0001101011111010",2374 => "0001101011111110",
2375 => "0001100001001101",2376 => "0001101100000101",
2377 => "0001101100001001",2378 => "0001101100001101",
2379 => "0001101100010001",2380 => "0001101100010101",
2381 => "0001101100011000",2382 => "0001101100011100",
2383 => "0001100000001000",2384 => "0001101100100100",
2385 => "0001101100101000",2386 => "0001101100101011",
2387 => "0001101100101111",2388 => "0001101100110011",
2389 => "0001101100110111",2390 => "0001101100111011",
2391 => "0001101100111111",2392 => "0001101101000010",
2393 => "0001101101000110",2394 => "0001101101001010",
2395 => "0001101101001110",2396 => "0001100001010101",
2397 => "0001101101010110",2398 => "0001101101011001",
2399 => "0001101101011101",2400 => "0001101101100001",
2401 => "0001101101100101",2402 => "0001101101101001",
2403 => "0001101101101101",2404 => "0001101101110001",
2405 => "0001101101110101",2406 => "0001101101111000",
2407 => "0001101101111100",2408 => "0001101110000000",
2409 => "0001100000001001",2410 => "0001101110001000",
2411 => "0001101110001100",2412 => "0001101110010000",
2413 => "0001101110010100",2414 => "0001100001011100",
2415 => "0001101110011100",2416 => "0001101110011111",
2417 => "0001101110100011",2418 => "0001101110100111",
2419 => "0001101110101011",2420 => "0001101110101111",
2421 => "0001101110110011",2422 => "0001101110110111",
2423 => "0001101110111011",2424 => "0001101110111111",
2425 => "0001101111000011",2426 => "0001101111000111",
2427 => "0001101111001011",2428 => "0001101111001111",
2429 => "0001101111010011",2430 => "0001101111010111",
2431 => "0001101111011011",2432 => "0001101111011111",
2433 => "0001101111100011",2434 => "0001101111100111",
2435 => "0010000000000011",2436 => "0010000000000111",
2437 => "0010000000001011",2438 => "0010000000001111",
2439 => "0010000000010011",2440 => "0010000000010111",
2441 => "0010000000011011",2442 => "0010000000011111",
2443 => "0010000000100011",2444 => "0010000000100111",
2445 => "0010000000101011",2446 => "0010000000101111",
2447 => "0010000000110011",2448 => "0010000000110111",
2449 => "0010000000111011",2450 => "0010000000111111",
2451 => "0010000001000011",2452 => "0010000001000111",
2453 => "0010000001001100",2454 => "0010000000001000",
2455 => "0010000001010100",2456 => "0010000001011000",
2457 => "0010000001011100",2458 => "0010000001100000",
2459 => "0010000000000001",2460 => "0010000001101000",
2461 => "0010000001101100",2462 => "0010000001110000",
2463 => "0010000001110100",2464 => "0010000001111001",
2465 => "0010000001111101",2466 => "0010000010000001",
2467 => "0010000010000101",2468 => "0010000010001001",
2469 => "0010000010001101",2470 => "0010000010010001",
2471 => "0010000000001111",2472 => "0010000010011010",
2473 => "0010000010011110",2474 => "0010000010100010",
2475 => "0010000010100110",2476 => "0010000000010001",
2477 => "0010000010101111",2478 => "0010000010110011",
2479 => "0010000010110111",2480 => "0010000010111011",
2481 => "0010000010111111",2482 => "0010000011000011",
2483 => "0010000000000010",2484 => "0010000011001100",
2485 => "0010000011010000",2486 => "0010000011010100",
2487 => "0010000011011000",2488 => "0010000011011101",
2489 => "0010000011100001",2490 => "0010000011100101",
2491 => "0010000011101001",2492 => "0010000011101110",
2493 => "0010000011110010",2494 => "0010000011110110",
2495 => "0010000000011001",2496 => "0010000011111111",
2497 => "0010000100000011",2498 => "0010000100000111",
2499 => "0010000100001011",2500 => "0010000100010000",
2501 => "0010000100010100",2502 => "0010000000011100",
2503 => "0010000100011100",2504 => "0010000100100001",
2505 => "0010000100100101",2506 => "0010000100101001",
2507 => "0010000100101110",2508 => "0010000100110010",
2509 => "0010000000011111",2510 => "0010000100111011",
2511 => "0010000100111111",2512 => "0010000101000011",
2513 => "0010000101001000",2514 => "0010000101001100",
2515 => "0010000101010000",2516 => "0010000101010101",
2517 => "0010000101011001",2518 => "0010000101011101",
2519 => "0010000101100010",2520 => "0010000101100110",
2521 => "0010000101101010",2522 => "0010000101101111",
2523 => "0010000101110011",2524 => "0010000101110111",
2525 => "0010000000100110",2526 => "0010000110000000",
2527 => "0010000110000101",2528 => "0010000110001001",
2529 => "0010000110001101",2530 => "0010000110010010",
2531 => "0010000110010110",2532 => "0010000110011011",
2533 => "0010000110011111",2534 => "0010000110100011",
2535 => "0010000110101000",2536 => "0010000110101100",
2537 => "0010000110110001",2538 => "0010000110110101",
2539 => "0010000110111010",2540 => "0010000110111110",
2541 => "0010000000101101",2542 => "0010000111000111",
2543 => "0010000111001011",2544 => "0010000111010000",
2545 => "0010000111010100",2546 => "0010000111011001",
2547 => "0010000111011101",2548 => "0010000111100010",
2549 => "0010000111100110",2550 => "0010000111101011",
2551 => "0010000111101111",2552 => "0010000000000101",
2553 => "0010000111111000",2554 => "0010000111111101",
2555 => "0010001000000001",2556 => "0010001000000110",
2557 => "0010001000001010",2558 => "0010001000001111",
2559 => "0010001000010011",2560 => "0010001000011000",
2561 => "0010000000110110",2562 => "0010001000100001",
2563 => "0010001000100101",2564 => "0010001000101010",
2565 => "0010001000101111",2566 => "0010001000110011",
2567 => "0010001000111000",2568 => "0010001000111100",
2569 => "0010001001000001",2570 => "0010001001000101",
2571 => "0010001001001010",2572 => "0010001001001111",
2573 => "0010001001010011",2574 => "0010000000000110",
2575 => "0010001001011100",2576 => "0010001001100001",
2577 => "0010001001100110",2578 => "0010001001101010",
2579 => "0010001001101111",2580 => "0010001001110011",
2581 => "0010001001111000",2582 => "0010001001111101",
2583 => "0010001010000001",2584 => "0010001010000110",
2585 => "0010001010001011",2586 => "0010001010001111",
2587 => "0010000001000010",2588 => "0010001010011001",
2589 => "0010001010011101",2590 => "0010001010100010",
2591 => "0010001010100111",2592 => "0010001010101011",
2593 => "0010001010110000",2594 => "0010001010110101",
2595 => "0010001010111001",2596 => "0010001010111110",
2597 => "0010001011000011",2598 => "0010001011000111",
2599 => "0010001011001100",2600 => "0010001011010001",
2601 => "0010001011010110",2602 => "0010000001001001",
2603 => "0010001011011111",2604 => "0010000001001010",
2605 => "0010001011101001",2606 => "0010001011101101",
2607 => "0010001011110010",2608 => "0010001011110111",
2609 => "0010001011111100",2610 => "0010001100000000",
2611 => "0010001100000101",2612 => "0010001100001010",
2613 => "0010001100001111",2614 => "0010001100010011",
2615 => "0010001100011000",2616 => "0010001100011101",
2617 => "0010001100100010",2618 => "0010001100100111",
2619 => "0010001100101011",2620 => "0010001100110000",
2621 => "0010001100110101",2622 => "0010001100111010",
2623 => "0010001100111111",2624 => "0010001101000100",
2625 => "0010000001010100",2626 => "0010001101001101",
2627 => "0010000001010101",2628 => "0010001101010111",
2629 => "0010000001010110",2630 => "0010001101100001",
2631 => "0010000001010111",2632 => "0010001101101010",
2633 => "0010001101101111",2634 => "0010001101110100",
2635 => "0010001101111001",2636 => "0010001101111110",
2637 => "0010001110000011",2638 => "0010001110001000",
2639 => "0010001110001101",2640 => "0010001110010010",
2641 => "0010001110010110",2642 => "0010001110011011",
2643 => "0010001110100000",2644 => "0010001110100101",
2645 => "0010001110101010",2646 => "0010001110101111",
2647 => "0010001110110100",2648 => "0010001110111001",
2649 => "0010001110111110",2650 => "0010001111000011",
2651 => "0010001111001000",2652 => "0010001111001101",
2653 => "0010001111010010",2654 => "0010001111010111",
2655 => "0010001111011100",2656 => "0010001111100001",
2657 => "0010001111100110",2658 => "0010100000000011",
2659 => "0010100000001000",2660 => "0010100000001101",
2661 => "0010100000010010",2662 => "0010100000010111",
2663 => "0010100000011100",2664 => "0010100000100001",
2665 => "0010100000100110",2666 => "0010100000101011",
2667 => "0010100000110000",2668 => "0010100000110101",
2669 => "0010100000111010",2670 => "0010100000111111",
2671 => "0010100001000100",2672 => "0010100001001001",
2673 => "0010100001001110",2674 => "0010100001010011",
2675 => "0010100001011001",2676 => "0010100001011110",
2677 => "0010100001100011",2678 => "0010100001101000",
2679 => "0010100001101101",2680 => "0010100001110010",
2681 => "0010100001110111",2682 => "0010100001111100",
2683 => "0010100010000001",2684 => "0010100010000111",
2685 => "0010100000001110",2686 => "0010100010010001",
2687 => "0010100000001111",2688 => "0010100010011011",
2689 => "0010100000010000",2690 => "0010100010100101",
2691 => "0010100010101011",2692 => "0010100010110000",
2693 => "0010100010110101",2694 => "0010100010111010",
2695 => "0010100010111111",2696 => "0010100011000101",
2697 => "0010100011001010",2698 => "0010100011001111",
2699 => "0010100011010100",2700 => "0010100011011001",
2701 => "0010100011011111",2702 => "0010100011100100",
2703 => "0010100011101001",2704 => "0010100011101110",
2705 => "0010100011110100",2706 => "0010100011111001",
2707 => "0010100011111110",2708 => "0010100100000011",
2709 => "0010100100001001",2710 => "0010100000011011",
2711 => "0010100100010011",2712 => "0010100000011100",
2713 => "0010100100011110",2714 => "0010100100100011",
2715 => "0010100100101000",2716 => "0010100100101110",
2717 => "0010100100110011",2718 => "0010100100111000",
2719 => "0010100100111101",2720 => "0010100101000011",
2721 => "0010100101001000",2722 => "0010100101001101",
2723 => "0010100101010011",2724 => "0010100101011000",
2725 => "0010100101011101",2726 => "0010100101100011",
2727 => "0010100000100100",2728 => "0010100101101110",
2729 => "0010100101110011",2730 => "0010100101111000",
2731 => "0010100101111110",2732 => "0010100110000011",
2733 => "0010100110001000",2734 => "0010100110001110",
2735 => "0010100110010011",2736 => "0010100110011001",
2737 => "0010100110011110",2738 => "0010100110100011",
2739 => "0010100110101001",2740 => "0010100000101011",
2741 => "0010100110110100",2742 => "0010100110111001",
2743 => "0010100110111111",2744 => "0010100111000100",
2745 => "0010100111001010",2746 => "0010100111001111",
2747 => "0010100111010100",2748 => "0010100111011010",
2749 => "0010100111011111",2750 => "0010100111100101",
2751 => "0010100000110001",2752 => "0010100111110000",
2753 => "0010100111110101",2754 => "0010100111111011",
2755 => "0010101000000000",2756 => "0010101000000110",
2757 => "0010101000001011",2758 => "0010101000010001",
2759 => "0010101000010110",2760 => "0010100000110110",
2761 => "0010101000100010",2762 => "0010101000100111",
2763 => "0010101000101101",2764 => "0010101000110010",
2765 => "0010101000111000",2766 => "0010101000111101",
2767 => "0010101001000011",2768 => "0010101001001001",
2769 => "0010100000111011",2770 => "0010101001010100",
2771 => "0010101001011001",2772 => "0010101001011111",
2773 => "0010101001100101",2774 => "0010101001101010",
2775 => "0010101001110000",2776 => "0010101001110101",
2777 => "0010101001111011",2778 => "0010101010000001",
2779 => "0010101010000110",2780 => "0010101010001100",
2781 => "0010101010010010",2782 => "0010101010010111",
2783 => "0010101010011101",2784 => "0010101010100011",
2785 => "0010100001000100",2786 => "0010101010101110",
2787 => "0010101010110100",2788 => "0010101010111001",
2789 => "0010101010111111",2790 => "0010101011000101",
2791 => "0010101011001010",2792 => "0010100001001000",
2793 => "0010101011010110",2794 => "0010101011011100",
2795 => "0010101011100001",2796 => "0010101011100111",
2797 => "0010101011101101",2798 => "0010101011110011",
2799 => "0010100001001100",2800 => "0010101011111110",
2801 => "0010101100000100",2802 => "0010101100001010",
2803 => "0010101100001111",2804 => "0010101100010101",
2805 => "0010101100011011",2806 => "0010101100100001",
2807 => "0010101100100111",2808 => "0010101100101100",
2809 => "0010101100110010",2810 => "0010101100111000",
2811 => "0010100001010011",2812 => "0010101101000100",
2813 => "0010101101001010",2814 => "0010101101001111",
2815 => "0010101101010101",2816 => "0010101101011011",
2817 => "0010101101100001",2818 => "0010101101100111",
2819 => "0010101101101101",2820 => "0010101101110011",
2821 => "0010101101111000",2822 => "0010101101111110",
2823 => "0010100000001001",2824 => "0010101110001010",
2825 => "0010101110010000",2826 => "0010101110010110",
2827 => "0010101110011100",2828 => "0010100001011101",
2829 => "0010101110101000",2830 => "0010101110101110",
2831 => "0010101110110100",2832 => "0010101110111010",
2833 => "0010100001100000",2834 => "0010101111000110",
2835 => "0010101111001100",2836 => "0010101111010001",
2837 => "0010101111010111",2838 => "0010101111011101",
2839 => "0010101111100011",2840 => "0011000000000001",
2841 => "0011000000000111",2842 => "0011000000001101",
2843 => "0011000000010011",2844 => "0011000000011001",
2845 => "0011000000100000",2846 => "0011000000100110",
2847 => "0011000000101100",2848 => "0011000000000101",
2849 => "0011000000111000",2850 => "0011000000111110",
2851 => "0011000001000100",2852 => "0011000001001010",
2853 => "0011000000001000",2854 => "0011000001010110",
2855 => "0011000001011100",2856 => "0011000001100010",
2857 => "0011000001101000",2858 => "0011000000001011",
2859 => "0011000001110101",2860 => "0011000001111011",
2861 => "0011000010000001",2862 => "0011000010000111",
2863 => "0011000010001101",2864 => "0011000010010011",
2865 => "0011000010011001",2866 => "0011000000010000",
2867 => "0011000010100110",2868 => "0011000010101100",
2869 => "0011000010110010",2870 => "0011000010111000",
2871 => "0011000000010011",2872 => "0011000011000101",
2873 => "0011000011001011",2874 => "0011000011010001",
2875 => "0011000011010111",2876 => "0011000011011101",
2877 => "0011000011100100",2878 => "0011000011101010",
2879 => "0011000000011000",2880 => "0011000011110110",
2881 => "0011000011111101",2882 => "0011000100000011",
2883 => "0011000100001001",2884 => "0011000100001111",
2885 => "0011000100010110",2886 => "0011000100011100",
2887 => "0011000000011101",2888 => "0011000100101001",
2889 => "0011000100101111",2890 => "0011000100110101",
2891 => "0011000100111011",2892 => "0011000101000010",
2893 => "0011000101001000",2894 => "0011000101001110",
2895 => "0011000101010101",2896 => "0011000101011011",
2897 => "0011000101100001",2898 => "0011000000100100",
2899 => "0011000101101110",2900 => "0011000101110101",
2901 => "0011000101111011",2902 => "0011000110000001",
2903 => "0011000110001000",2904 => "0011000110001110",
2905 => "0011000110010100",2906 => "0011000110011011",
2907 => "0011000110100001",2908 => "0011000110101000",
2909 => "0011000000101011",2910 => "0011000110110101",
2911 => "0011000110111011",2912 => "0011000111000001",
2913 => "0011000111001000",2914 => "0011000111001110",
2915 => "0011000111010101",2916 => "0011000111011011",
2917 => "0011000111100010",2918 => "0011000111101000",
2919 => "0011000111101111",2920 => "0011000111110101",
2921 => "0011000111111100",2922 => "0011001000000010",
2923 => "0011001000001001",2924 => "0011001000001111",
2925 => "0011001000010110",2926 => "0011000000110110",
2927 => "0011001000100011",2928 => "0011001000101010",
2929 => "0011000000111000",2930 => "0011001000110111",
2931 => "0011001000111101",2932 => "0011000000111010",
2933 => "0011001001001010",2934 => "0011001001010001",
2935 => "0011000000000110",2936 => "0011001001011110",
2937 => "0011001001100101",2938 => "0011001001101011",
2939 => "0011001001110010",2940 => "0011001001111001",
2941 => "0011001001111111",2942 => "0011001010000110",
2943 => "0011001010001101",2944 => "0011001010010011",
2945 => "0011001010011010",2946 => "0011001010100001",
2947 => "0011001010100111",2948 => "0011001010101110",
2949 => "0011001010110101",2950 => "0011001010111011",
2951 => "0011001011000010",2952 => "0011001011001001",
2953 => "0011001011001111",2954 => "0011001011010110",
2955 => "0011001011011101",2956 => "0011000001001010",
2957 => "0011001011101010",2958 => "0011001011110001",
2959 => "0011000001001100",2960 => "0011001011111111",
2961 => "0011001100000101",2962 => "0011000001001110",
2963 => "0011001100010011",2964 => "0011001100011010",
2965 => "0011001100100001",2966 => "0011001100100111",
2967 => "0011001100101110",2968 => "0011001100110101",
2969 => "0011001100111100",2970 => "0011001101000011",
2971 => "0011001101001001",2972 => "0011001101010000",
2973 => "0011001101010111",2974 => "0011001101011110",
2975 => "0011001101100101",2976 => "0011001101101100",
2977 => "0011001101110011",2978 => "0011000001011001",
2979 => "0011001110000000",2980 => "0011001110000111",
2981 => "0011000001011011",2982 => "0011001110010101",
2983 => "0011001110011100",2984 => "0011001110100011",
2985 => "0011001110101010",2986 => "0011001110110001",
2987 => "0011001110111000",2988 => "0011001110111111",
2989 => "0011001111000110",2990 => "0011001111001101",
2991 => "0011000001100010",2992 => "0011001111011011",
2993 => "0011001111100010",2994 => "0011100000000001",
2995 => "0011100000001000",2996 => "0011100000001111",
2997 => "0011100000010110",2998 => "0011100000011101",
2999 => "0011100000100100",3000 => "0011100000101011",
3001 => "0011100000000101",3002 => "0011100000111001",
3003 => "0011100001000000",3004 => "0011100001000111",
3005 => "0011100001001110",3006 => "0011100001010101",
3007 => "0011100001011100",3008 => "0011100001100011",
3009 => "0011100001101010",3010 => "0011100001110010",
3011 => "0011100001111001",3012 => "0011100010000000",
3013 => "0011100010000111",3014 => "0011100010001110",
3015 => "0011100010010101",3016 => "0011100010011100",
3017 => "0011100010100100",3018 => "0011100010101011",
3019 => "0011100010110010",3020 => "0011100010111001",
3021 => "0011100011000000",3022 => "0011100011000111",
3023 => "0011100011001111",3024 => "0011100011010110",
3025 => "0011100011011101",3026 => "0011100011100100",
3027 => "0011100011101100",3028 => "0011100011110011",
3029 => "0011100000011001",3030 => "0011100100000001",
3031 => "0011100100001001",3032 => "0011100100010000",
3033 => "0011100100010111",3034 => "0011100100011110",
3035 => "0011100100100110",3036 => "0011100100101101",
3037 => "0011100100110100",3038 => "0011100100111100",
3039 => "0011100101000011",3040 => "0011100000100001",
3041 => "0011100101010010",3042 => "0011100101011001",
3043 => "0011100101100000",3044 => "0011100000100100",
3045 => "0011100101101111",3046 => "0011100101110110",
3047 => "0011100101111110",3048 => "0001100000000100",
3049 => "0001100000000100",3050 => "0001100000000101",
3051 => "0001100000000101",3052 => "0001100000000101",
3053 => "0001100000000110",3054 => "0001100000000110",
3055 => "0001100000000110",3056 => "0001100000000111",
3057 => "0001100000000111",3058 => "0001100000000111",
3059 => "0001100000000111",3060 => "0001100000001000",
3061 => "0001100000001000",3062 => "0001100000001000",
3063 => "0001100000001001",3064 => "0001100000001001",
3065 => "0001100000001001",3066 => "0001100000000001",
3067 => "0001100000000001",3068 => "0001100000000001",
3069 => "0001100000000001",3070 => "0001100000001011",
3071 => "0001100000001011",3072 => "0001100000001011",
3073 => "0001100000001100",3074 => "0001100000001100",
3075 => "0001100000001100",3076 => "0001100000001101",
3077 => "0001100000001101",3078 => "0001100000001101",
3079 => "0001100000001101",3080 => "0001100000001110",
3081 => "0001100000001110",3082 => "0001100000001110",
3083 => "0001100000001111",3084 => "0001100000001111",
3085 => "0001100000001111",3086 => "0001100000010000",
3087 => "0001100000010000",3088 => "0001100000010000",
3089 => "0001100000010001",3090 => "0001100000010001",
3091 => "0001100000010001",3092 => "0001100000010001",
3093 => "0001100000010010",3094 => "0001100000010010",
3095 => "0001100000010010",3096 => "0001100000010011",
3097 => "0001100000010011",3098 => "0001100000010011",
3099 => "0001100000000010",3100 => "0001100000000010",
3101 => "0001100000000010",3102 => "0001100000000010",
3103 => "0001100000010101",3104 => "0001100000010101",
3105 => "0001100000010101",3106 => "0001100000010110",
3107 => "0001100000010110",3108 => "0001100000010110",
3109 => "0001100000010111",3110 => "0001100000010111",
3111 => "0001100000010111",3112 => "0001100000010111",
3113 => "0001100000011000",3114 => "0001100000011000",
3115 => "0001100000011000",3116 => "0001100000011001",
3117 => "0001100000011001",3118 => "0001100000011001",
3119 => "0001100000011010",3120 => "0001100000011010",
3121 => "0001100000011010",3122 => "0001100000011010",
3123 => "0001100000011011",3124 => "0001100000011011",
3125 => "0001100000011011",3126 => "0001100000011100",
3127 => "0001100000011100",3128 => "0001100000011100",
3129 => "0001100000011101",3130 => "0001100000011101",
3131 => "0001100000011101",3132 => "0001100000000011",
3133 => "0001100000000011",3134 => "0001100000000011",
3135 => "0001100000000011",3136 => "0001100000011111",
3137 => "0001100000011111",3138 => "0001100000011111",
3139 => "0001100000100000",3140 => "0001100000100000",
3141 => "0001100000100000",3142 => "0001100000100001",
3143 => "0001100000100001",3144 => "0001100000100001",
3145 => "0001100000100001",3146 => "0001100000100010",
3147 => "0001100000100010",3148 => "0001100000100010",
3149 => "0001100000100011",3150 => "0001100000100011",
3151 => "0001100000100011",3152 => "0001100000100100",
3153 => "0001100000100100",3154 => "0001100000100100",
3155 => "0001100000100100",3156 => "0001100000100101",
3157 => "0001100000100101",3158 => "0001100000100101",
3159 => "0001100000100110",3160 => "0001100000100110",
3161 => "0001100000100110",3162 => "0001100000100111",
3163 => "0001100000100111",3164 => "0001100000100111",
3165 => "0001100000000100",3166 => "0001100000000100",
3167 => "0001100000000100",3168 => "0001100000000100",
3169 => "0001100000101001",3170 => "0001100000101001",
3171 => "0001100000101001",3172 => "0001100000101010",
3173 => "0001100000101010",3174 => "0001100000101010",
3175 => "0001100000101011",3176 => "0001100000101011",
3177 => "0001100000101011",3178 => "0001100000101011",
3179 => "0001100000101100",3180 => "0001100000101100",
3181 => "0001100000101100",3182 => "0001100000101101",
3183 => "0001100000101101",3184 => "0001100000101101",
3185 => "0001100000101110",3186 => "0001100000101110",
3187 => "0001100000101110",3188 => "0001100000101111",
3189 => "0001100000101111",3190 => "0001100000101111",
3191 => "0001100000101111",3192 => "0001100000110000",
3193 => "0001100000110000",3194 => "0001100000110000",
3195 => "0001100000110001",3196 => "0001100000110001",
3197 => "0001100000110001",3198 => "0001100000000101",
3199 => "0001100000000101",3200 => "0001100000000101",
3201 => "0001100000000101",3202 => "0001100000110011",
3203 => "0001100000110011",3204 => "0001100000110011",
3205 => "0001100000110100",3206 => "0001100000110100",
3207 => "0001100000110100",3208 => "0001100000110101",
3209 => "0001100000110101",3210 => "0001100000110101",
3211 => "0001100000110110",3212 => "0001100000110110",
3213 => "0001100000110110",3214 => "0001100000110110",
3215 => "0001100000110111",3216 => "0001100000110111",
3217 => "0001100000110111",3218 => "0001100000111000",
3219 => "0001100000111000",3220 => "0001100000111000",
3221 => "0001100000111001",3222 => "0001100000111001",
3223 => "0001100000111001",3224 => "0001100000111010",
3225 => "0001100000111010",3226 => "0001100000111010",
3227 => "0001100000111010",3228 => "0001100000111011",
3229 => "0001100000111011",3230 => "0001100000111011",
3231 => "0001100000000110",3232 => "0001100000000110",
3233 => "0001100000000110",3234 => "0001100000111101",
3235 => "0001100000111101",3236 => "0001100000111101",
3237 => "0001100000111101",3238 => "0001100000111110",
3239 => "0001100000111110",3240 => "0001100000111110",
3241 => "0001100000111111",3242 => "0001100000111111",
3243 => "0001100000111111",3244 => "0001100001000000",
3245 => "0001100001000000",3246 => "0001100001000000",
3247 => "0001100001000001",3248 => "0001100001000001",
3249 => "0001100001000001",3250 => "0001100001000001",
3251 => "0001100001000010",3252 => "0001100001000010",
3253 => "0001100001000010",3254 => "0001100001000011",
3255 => "0001100001000011",3256 => "0001100001000011",
3257 => "0001100001000100",3258 => "0001100001000100",
3259 => "0001100001000100",3260 => "0001100001000101",
3261 => "0001100001000101",3262 => "0001100001000101",
3263 => "0001100001000101",3264 => "0001100000000111",
3265 => "0001100000000111",3266 => "0001100000000111",
3267 => "0001100001000111",3268 => "0001100001000111",
3269 => "0001100001000111",3270 => "0001100001001000",
3271 => "0001100001001000",3272 => "0001100001001000",
3273 => "0001100001001001",3274 => "0001100001001001",
3275 => "0001100001001001",3276 => "0001100001001001",
3277 => "0001100001001010",3278 => "0001100001001010",
3279 => "0001100001001010",3280 => "0001100001001011",
3281 => "0001100001001011",3282 => "0001100001001011",
3283 => "0001100001001100",3284 => "0001100001001100",
3285 => "0001100001001100",3286 => "0001100001001101",
3287 => "0001100001001101",3288 => "0001100001001101",
3289 => "0001100001001101",3290 => "0001100001001110",
3291 => "0001100001001110",3292 => "0001100001001110",
3293 => "0001100001001111",3294 => "0001100001001111",
3295 => "0001100001001111",3296 => "0001100000001000",
3297 => "0001100000001000",3298 => "0001100000001000",
3299 => "0001100001010001",3300 => "0001100001010001",
3301 => "0001100001010001",3302 => "0001100001010001",
3303 => "0001100001010010",3304 => "0001100001010010",
3305 => "0001100001010010",3306 => "0001100001010011",
3307 => "0001100001010011",3308 => "0001100001010011",
3309 => "0001100001010100",3310 => "0001100001010100",
3311 => "0001100001010100",3312 => "0001100001010101",
3313 => "0001100001010101",3314 => "0001100001010101",
3315 => "0001100001010101",3316 => "0001100001010110",
3317 => "0001100001010110",3318 => "0001100001010110",
3319 => "0001100001010111",3320 => "0001100001010111",
3321 => "0001100001010111",3322 => "0001100001011000",
3323 => "0001100001011000",3324 => "0001100001011000",
3325 => "0001100001011001",3326 => "0001100001011001",
3327 => "0001100001011001",3328 => "0001100001011001",
3329 => "0001100000001001",3330 => "0001100000001001",
3331 => "0001100000001001",3332 => "0001100001011011",
3333 => "0001100001011011",3334 => "0001100001011011",
3335 => "0001100001011100",3336 => "0001100001011100",
3337 => "0001100001011100",3338 => "0001100001011101",
3339 => "0001100001011101",3340 => "0001100001011101",
3341 => "0001100001011101",3342 => "0001100001011110",
3343 => "0001100001011110",3344 => "0001100001011110",
3345 => "0001100001011111",3346 => "0001100001011111",
3347 => "0001100001011111",3348 => "0001100001100000",
3349 => "0001100001100000",3350 => "0001100001100000",
3351 => "0001100001100001",3352 => "0001100001100001",
3353 => "0001100001100001",3354 => "0001100001100010",
3355 => "0001100001100010",3356 => "0001100001100010",
3357 => "0001100001100010",3358 => "0001100001100011",
3359 => "0001100001100011",3360 => "0001100001100011",
3361 => "0001100000000001",3362 => "0001100000000001",
3363 => "0001100000000001",3364 => "0001100001100101",
3365 => "0001100001100101",3366 => "0001100001100101",
3367 => "0001100001100110",3368 => "0001100001100110",
3369 => "0001100001100110",3370 => "0001100001100110",
3371 => "0001100001100111",3372 => "0001100001100111",
3373 => "0001100001100111",3374 => "0001100001101000",
3375 => "0001100001101000",3376 => "0001100001101000",
3377 => "0001100001101001",3378 => "0001100001101001",
3379 => "0001100001101001",3380 => "0001100001101010",
3381 => "0001100001101010",3382 => "0001100001101010",
3383 => "0001100001101011",3384 => "0001100001101011",
3385 => "0001100001101011",3386 => "0001100001101011",
3387 => "0001100001101100",3388 => "0001100001101100",
3389 => "0001100001101100",3390 => "0001100001101101",
3391 => "0001100001101101",3392 => "0001100001101101",
3393 => "0001100000001011",3394 => "0001100000001011",
3395 => "0001100000001011",3396 => "0001100001101111",
3397 => "0001100001101111",3398 => "0001100001101111",
3399 => "0001100001101111",3400 => "0001100001110000",
3401 => "0001100001110000",3402 => "0001100001110000",
3403 => "0001100001110001",3404 => "0001100001110001",
3405 => "0001100001110001",3406 => "0001100001110010",
3407 => "0001100001110010",3408 => "0001100001110010",
3409 => "0001100001110011",3410 => "0001100001110011",
3411 => "0001100001110011",3412 => "0001100001110100",
3413 => "0001100001110100",3414 => "0001100001110100",
3415 => "0001100001110100",3416 => "0001100001110101",
3417 => "0001100001110101",3418 => "0001100001110101",
3419 => "0001100001110110",3420 => "0001100001110110",
3421 => "0001100001110110",3422 => "0001100001110111",
3423 => "0001100001110111",3424 => "0001100001110111",
3425 => "0001100000001100",3426 => "0001100000001100",
3427 => "0001100000001100",3428 => "0001100001111001",
3429 => "0001100001111001",3430 => "0001100001111001",
3431 => "0001100001111001",3432 => "0001100001111010",
3433 => "0001100001111010",3434 => "0001100001111010",
3435 => "0001100001111011",3436 => "0001100001111011",
3437 => "0001100001111011",3438 => "0001100001111100",
3439 => "0001100001111100",3440 => "0001100001111100",
3441 => "0001100001111101",3442 => "0001100001111101",
3443 => "0001100001111101",3444 => "0001100001111110",
3445 => "0001100001111110",3446 => "0001100001111110",
3447 => "0001100001111110",3448 => "0001100001111111",
3449 => "0001100001111111",3450 => "0001100001111111",
3451 => "0001100010000000",3452 => "0001100010000000",
3453 => "0001100010000000",3454 => "0001100010000001",
3455 => "0001100010000001",3456 => "0001100010000001",
3457 => "0001100000001101",3458 => "0001100000001101",
3459 => "0001100000001101",3460 => "0001100010000011",
3461 => "0001100010000011",3462 => "0001100010000011",
3463 => "0001100010000011",3464 => "0001100010000100",
3465 => "0001100010000100",3466 => "0001100010000100",
3467 => "0001100010000101",3468 => "0001100010000101",
3469 => "0001100010000101",3470 => "0001100010000110",
3471 => "0001100010000110",3472 => "0001100010000110",
3473 => "0001100010000111",3474 => "0001100010000111",
3475 => "0001100010000111",3476 => "0001100010001000",
3477 => "0001100010001000",3478 => "0001100010001000",
3479 => "0001100010001000",3480 => "0001100010001001",
3481 => "0001100010001001",3482 => "0001100010001001",
3483 => "0001100010001010",3484 => "0001100010001010",
3485 => "0001100010001010",3486 => "0001100010001011",
3487 => "0001100010001011",3488 => "0001100010001011",
3489 => "0001100000001110",3490 => "0001100000001110",
3491 => "0001100000001110",3492 => "0001100010001101",
3493 => "0001100010001101",3494 => "0001100010001101",
3495 => "0001100010001101",3496 => "0001100010001110",
3497 => "0001100010001110",3498 => "0001100010001110",
3499 => "0001100010001111",3500 => "0001100010001111",
3501 => "0001100010001111",3502 => "0001100010010000",
3503 => "0001100010010000",3504 => "0001100010010000",
3505 => "0001100010010001",3506 => "0001100010010001",
3507 => "0001100010010001",3508 => "0001100010010010",
3509 => "0001100010010010",3510 => "0001100010010010",
3511 => "0001100010010011",3512 => "0001100010010011",
3513 => "0001100010010011",3514 => "0001100010010011",
3515 => "0001100010010100",3516 => "0001100010010100",
3517 => "0001100010010100",3518 => "0001100010010101",
3519 => "0001100010010101",3520 => "0001100010010101",
3521 => "0001100000001111",3522 => "0001100000001111",
3523 => "0001100000001111",3524 => "0001100010010111",
3525 => "0001100010010111",3526 => "0001100010010111",
3527 => "0001100010011000",3528 => "0001100010011000",
3529 => "0001100010011000",3530 => "0001100010011001",
3531 => "0001100010011001",3532 => "0001100010011001",
3533 => "0001100010011001",3534 => "0001100010011010",
3535 => "0001100010011010",3536 => "0001100010011010",
3537 => "0001100010011011",3538 => "0001100010011011",
3539 => "0001100010011011",3540 => "0001100010011100",
3541 => "0001100010011100",3542 => "0001100010011100",
3543 => "0001100010011101",3544 => "0001100010011101",
3545 => "0001100010011101",3546 => "0001100010011110",
3547 => "0001100010011110",3548 => "0001100010011110",
3549 => "0001100010011111",3550 => "0001100010011111",
3551 => "0001100010011111",3552 => "0001100010011111",
3553 => "0001100000010000",3554 => "0001100000010000",
3555 => "0001100000010000",3556 => "0001100010100001",
3557 => "0001100010100001",3558 => "0001100010100001",
3559 => "0001100010100010",3560 => "0001100010100010",
3561 => "0001100010100010",3562 => "0001100010100011",
3563 => "0001100010100011",3564 => "0001100010100011",
3565 => "0001100010100100",3566 => "0001100010100100",
3567 => "0001100010100100",3568 => "0001100010100101",
3569 => "0001100010100101",3570 => "0001100010100101",
3571 => "0001100010100101",3572 => "0001100010100110",
3573 => "0001100010100110",3574 => "0001100010100110",
3575 => "0001100010100111",3576 => "0001100010100111",
3577 => "0001100010100111",3578 => "0001100010101000",
3579 => "0001100010101000",3580 => "0001100010101000",
3581 => "0001100010101001",3582 => "0001100010101001",
3583 => "0001100010101001",3584 => "0001100000010001",
3585 => "0001100000010001",3586 => "0001100000010001",
3587 => "0001100010101011",3588 => "0001100010101011",
3589 => "0001100010101011",3590 => "0001100010101011",
3591 => "0001100010101100",3592 => "0001100010101100",
3593 => "0001100010101100",3594 => "0001100010101101",
3595 => "0001100010101101",3596 => "0001100010101101",
3597 => "0001100010101110",3598 => "0001100010101110",
3599 => "0001100010101110",3600 => "0001100010101111",
3601 => "0001100010101111",3602 => "0001100010101111",
3603 => "0001100010110000",3604 => "0001100010110000",
3605 => "0001100010110000",3606 => "0001100010110001",
3607 => "0001100010110001",3608 => "0001100010110001",
3609 => "0001100010110010",3610 => "0001100010110010",
3611 => "0001100010110010",3612 => "0001100010110010",
3613 => "0001100010110011",3614 => "0001100010110011",
3615 => "0001100010110011",3616 => "0001100000010010",
3617 => "0001100000010010",3618 => "0001100000010010",
3619 => "0001100010110101",3620 => "0001100010110101",
3621 => "0001100010110101",3622 => "0001100010110110",
3623 => "0001100010110110",3624 => "0001100010110110",
3625 => "0001100010110111",3626 => "0001100010110111",
3627 => "0001100010110111",3628 => "0001100010111000",
3629 => "0001100010111000",3630 => "0001100010111000",
3631 => "0001100010111001",3632 => "0001100010111001",
3633 => "0001100010111001",3634 => "0001100010111001",
3635 => "0001100010111010",3636 => "0001100010111010",
3637 => "0001100010111010",3638 => "0001100010111011",
3639 => "0001100010111011",3640 => "0001100010111011",
3641 => "0001100010111100",3642 => "0001100010111100",
3643 => "0001100010111100",3644 => "0001100010111101",
3645 => "0001100010111101",3646 => "0001100010111101",
3647 => "0001100000010011",3648 => "0001100000010011",
3649 => "0001100000010011",3650 => "0001100010111111",
3651 => "0001100010111111",3652 => "0001100010111111",
3653 => "0001100011000000",3654 => "0001100011000000",
3655 => "0001100011000000",3656 => "0001100011000000",
3657 => "0001100011000001",3658 => "0001100011000001",
3659 => "0001100011000001",3660 => "0001100011000010",
3661 => "0001100011000010",3662 => "0001100011000010",
3663 => "0001100011000011",3664 => "0001100011000011",
3665 => "0001100011000011",3666 => "0001100011000100",
3667 => "0001100011000100",3668 => "0001100011000100",
3669 => "0001100011000101",3670 => "0001100011000101",
3671 => "0001100011000101",3672 => "0001100011000110",
3673 => "0001100011000110",3674 => "0001100011000110",
3675 => "0001100011000111",3676 => "0001100011000111",
3677 => "0001100011000111",3678 => "0001100000000010",
3679 => "0001100000000010",3680 => "0001100000000010",
3681 => "0001100000000010",3682 => "0001100011001001",
3683 => "0001100011001001",3684 => "0001100011001001",
3685 => "0001100011001010",3686 => "0001100011001010",
3687 => "0001100011001010",3688 => "0001100011001011",
3689 => "0001100011001011",3690 => "0001100011001011",
3691 => "0001100011001100",3692 => "0001100011001100",
3693 => "0001100011001100",3694 => "0001100011001101",
3695 => "0001100011001101",3696 => "0001100011001101",
3697 => "0001100011001110",3698 => "0001100011001110",
3699 => "0001100011001110",3700 => "0001100011001111",
3701 => "0001100011001111",3702 => "0001100011001111",
3703 => "0001100011010000",3704 => "0001100011010000",
3705 => "0001100011010000",3706 => "0001100011010000",
3707 => "0001100011010001",3708 => "0001100011010001",
3709 => "0001100011010001",3710 => "0001100000010101",
3711 => "0001100000010101",3712 => "0001100000010101",
3713 => "0001100011010011",3714 => "0001100011010011",
3715 => "0001100011010011",3716 => "0001100011010100",
3717 => "0001100011010100",3718 => "0001100011010100",
3719 => "0001100011010101",3720 => "0001100011010101",
3721 => "0001100011010101",3722 => "0001100011010110",
3723 => "0001100011010110",3724 => "0001100011010110",
3725 => "0001100011010111",3726 => "0001100011010111",
3727 => "0001100011010111",3728 => "0001100011011000",
3729 => "0001100011011000",3730 => "0001100011011000",
3731 => "0001100011011001",3732 => "0001100011011001",
3733 => "0001100011011001",3734 => "0001100011011001",
3735 => "0001100011011010",3736 => "0001100011011010",
3737 => "0001100011011010",3738 => "0001100011011011",
3739 => "0001100011011011",3740 => "0001100011011011",
3741 => "0001100000010110",3742 => "0001100000010110",
3743 => "0001100000010110",3744 => "0001100011011101",
3745 => "0001100011011101",3746 => "0001100011011101",
3747 => "0001100011011110",3748 => "0001100011011110",
3749 => "0001100011011110",3750 => "0001100011011111",
3751 => "0001100011011111",3752 => "0001100011011111",
3753 => "0001100011100000",3754 => "0001100011100000",
3755 => "0001100011100000",3756 => "0001100011100001",
3757 => "0001100011100001",3758 => "0001100011100001",
3759 => "0001100011100010",3760 => "0001100011100010",
3761 => "0001100011100010",3762 => "0001100011100011",
3763 => "0001100011100011",3764 => "0001100011100011",
3765 => "0001100011100011",3766 => "0001100011100100",
3767 => "0001100011100100",3768 => "0001100011100100",
3769 => "0001100011100101",3770 => "0001100011100101",
3771 => "0001100011100101",3772 => "0001100000010111",
3773 => "0001100000010111",3774 => "0001100000010111",
3775 => "0001100011100111",3776 => "0001100011100111",
3777 => "0001100011100111",3778 => "0001100011101000",
3779 => "0001100011101000",3780 => "0001100011101000",
3781 => "0001100011101001",3782 => "0001100011101001",
3783 => "0001100011101001",3784 => "0001100011101010",
3785 => "0001100011101010",3786 => "0001100011101010",
3787 => "0001100011101011",3788 => "0001100011101011",
3789 => "0001100011101011",3790 => "0001100011101100",
3791 => "0001100011101100",3792 => "0001100011101100",
3793 => "0001100011101101",3794 => "0001100011101101",
3795 => "0001100011101101",3796 => "0001100011101101",
3797 => "0001100011101110",3798 => "0001100011101110",
3799 => "0001100011101110",3800 => "0001100011101111",
3801 => "0001100011101111",3802 => "0001100011101111",
3803 => "0001100000011000",3804 => "0001100000011000",
3805 => "0001100000011000",3806 => "0001100011110001",
3807 => "0001100011110001",3808 => "0001100011110001",
3809 => "0001100011110010",3810 => "0001100011110010",
3811 => "0001100011110010",3812 => "0001100011110011",
3813 => "0001100011110011",3814 => "0001100011110011",
3815 => "0001100011110100",3816 => "0001100011110100",
3817 => "0001100011110100",3818 => "0001100011110101",
3819 => "0001100011110101",3820 => "0001100011110101",
3821 => "0001100011110110",3822 => "0001100011110110",
3823 => "0001100011110110",3824 => "0001100011110111",
3825 => "0001100011110111",3826 => "0001100011110111",
3827 => "0001100011111000",3828 => "0001100011111000",
3829 => "0001100011111000",3830 => "0001100011111001",
3831 => "0001100011111001",3832 => "0001100011111001",
3833 => "0001100011111001",3834 => "0001100000011001",
3835 => "0001100000011001",3836 => "0001100000011001",
3837 => "0001100011111011",3838 => "0001100011111011",
3839 => "0001100011111011",3840 => "0001100011111100",
3841 => "0001100011111100",3842 => "0001100011111100",
3843 => "0001100011111101",3844 => "0001100011111101",
3845 => "0001100011111101",3846 => "0001100011111110",
3847 => "0001100011111110",3848 => "0001100011111110",
3849 => "0001100011111111",3850 => "0001100011111111",
3851 => "0001100011111111",3852 => "0001100100000000",
3853 => "0001100100000000",3854 => "0001100100000000",
3855 => "0001100100000001",3856 => "0001100100000001",
3857 => "0001100100000001",3858 => "0001100100000010",
3859 => "0001100100000010",3860 => "0001100100000010",
3861 => "0001100100000011",3862 => "0001100100000011",
3863 => "0001100100000011",3864 => "0001100000011010",
3865 => "0001100000011010",3866 => "0001100000011010",
3867 => "0001100100000101",3868 => "0001100100000101",
3869 => "0001100100000101",3870 => "0001100100000110",
3871 => "0001100100000110",3872 => "0001100100000110",
3873 => "0001100100000111",3874 => "0001100100000111",
3875 => "0001100100000111",3876 => "0001100100000111",
3877 => "0001100100001000",3878 => "0001100100001000",
3879 => "0001100100001000",3880 => "0001100100001001",
3881 => "0001100100001001",3882 => "0001100100001001",
3883 => "0001100100001010",3884 => "0001100100001010",
3885 => "0001100100001010",3886 => "0001100100001011",
3887 => "0001100100001011",3888 => "0001100100001011",
3889 => "0001100100001100",3890 => "0001100100001100",
3891 => "0001100100001100",3892 => "0001100100001101",
3893 => "0001100100001101",3894 => "0001100100001101",
3895 => "0001100000011011",3896 => "0001100000011011",
3897 => "0001100000011011",3898 => "0001100100001111",
3899 => "0001100100001111",3900 => "0001100100001111",
3901 => "0001100100010000",3902 => "0001100100010000",
3903 => "0001100100010000",3904 => "0001100100010001",
3905 => "0001100100010001",3906 => "0001100100010001",
3907 => "0001100100010010",3908 => "0001100100010010",
3909 => "0001100100010010",3910 => "0001100100010011",
3911 => "0001100100010011",3912 => "0001100100010011",
3913 => "0001100100010100",3914 => "0001100100010100",
3915 => "0001100100010100",3916 => "0001100100010101",
3917 => "0001100100010101",3918 => "0001100100010101",
3919 => "0001100100010110",3920 => "0001100100010110",
3921 => "0001100100010110",3922 => "0001100100010111",
3923 => "0001100100010111",3924 => "0001100100010111",
3925 => "0001100000011100",3926 => "0001100000011100",
3927 => "0001100000011100",3928 => "0001100100011001",
3929 => "0001100100011001",3930 => "0001100100011001",
3931 => "0001100100011001",3932 => "0001100100011010",
3933 => "0001100100011010",3934 => "0001100100011010",
3935 => "0001100100011011",3936 => "0001100100011011",
3937 => "0001100100011011",3938 => "0001100100011100",
3939 => "0001100100011100",3940 => "0001100100011100",
3941 => "0001100100011101",3942 => "0001100100011101",
3943 => "0001100100011101",3944 => "0001100100011110",
3945 => "0001100100011110",3946 => "0001100100011110",
3947 => "0001100100011111",3948 => "0001100100011111",
3949 => "0001100100011111",3950 => "0001100100100000",
3951 => "0001100100100000",3952 => "0001100100100000",
3953 => "0001100100100001",3954 => "0001100100100001",
3955 => "0001100100100001",3956 => "0001100000011101",
3957 => "0001100000011101",3958 => "0001100000011101",
3959 => "0001100100100011",3960 => "0001100100100011",
3961 => "0001100100100011",3962 => "0001100100100100",
3963 => "0001100100100100",3964 => "0001100100100100",
3965 => "0001100100100101",3966 => "0001100100100101",
3967 => "0001100100100101",3968 => "0001100100100110",
3969 => "0001100100100110",3970 => "0001100100100110",
3971 => "0001100100100111",3972 => "0001100100100111",
3973 => "0001100100100111",3974 => "0001100100101000",
3975 => "0001100100101000",3976 => "0001100100101000",
3977 => "0001100100101001",3978 => "0001100100101001",
3979 => "0001100100101001",3980 => "0001100100101010",
3981 => "0001100100101010",3982 => "0001100100101010",
3983 => "0001100100101011",3984 => "0001100100101011",
3985 => "0001100100101011",3986 => "0001100000000011",
3987 => "0001100000000011",3988 => "0001100000000011",
3989 => "0001100100101101",3990 => "0001100100101101",
3991 => "0001100100101101",3992 => "0001100100101110",
3993 => "0001100100101110",3994 => "0001100100101110",
3995 => "0001100100101111",3996 => "0001100100101111",
3997 => "0001100100101111",3998 => "0001100100110000",
3999 => "0001100100110000",4000 => "0001100100110000",
4001 => "0001100100110001",4002 => "0001100100110001",
4003 => "0001100100110001",4004 => "0001100100110010",
4005 => "0001100100110010",4006 => "0001100100110010",
4007 => "0001100100110011",4008 => "0001100100110011",
4009 => "0001100100110011",4010 => "0001100100110100",
4011 => "0001100100110100",4012 => "0001100100110100",
4013 => "0001100100110101",4014 => "0001100100110101",
4015 => "0001100100110101",4016 => "0001100000011111",
4017 => "0001100000011111",4018 => "0001100000011111",
4019 => "0001100100110111",4020 => "0001100100110111",
4021 => "0001100100110111",4022 => "0001100100110111",
4023 => "0001100100111000",4024 => "0001100100111000",
4025 => "0001100100111000",4026 => "0001100100111001",
4027 => "0001100100111001",4028 => "0001100100111001",
4029 => "0001100100111010",4030 => "0001100100111010",
4031 => "0001100100111010",4032 => "0001100100111011",
4033 => "0001100100111011",4034 => "0001100100111011",
4035 => "0001100100111100",4036 => "0001100100111100",
4037 => "0001100100111100",4038 => "0001100100111101",
4039 => "0001100100111101",4040 => "0001100100111101",
4041 => "0001100100111110",4042 => "0001100100111110",
4043 => "0001100100111110",4044 => "0001100100111111",
4045 => "0001100100111111",4046 => "0001100100111111",
4047 => "0001100000100000",4048 => "0001100000100000",
4049 => "0001100000100000",4050 => "0001100101000001",
4051 => "0001100101000001",4052 => "0001100101000001",
4053 => "0001100101000010",4054 => "0001100101000010",
4055 => "0001100101000010",4056 => "0001100101000011",
4057 => "0001100101000011",4058 => "0001100101000011",
4059 => "0001100101000100",4060 => "0001100101000100",
4061 => "0001100101000100",4062 => "0001100101000101",
4063 => "0001100101000101",4064 => "0001100101000101",
4065 => "0001100101000110",4066 => "0001100101000110",
4067 => "0001100101000110",4068 => "0001100101000111",
4069 => "0001100101000111",4070 => "0001100101000111",
4071 => "0001100101001000",4072 => "0001100101001000",
4073 => "0001100101001000",4074 => "0001100101001001",
4075 => "0001100101001001",4076 => "0001100101001001",
4077 => "0001100000100001",4078 => "0001100000100001",
4079 => "0001100000100001",4080 => "0001100101001011",
4081 => "0001100101001011",4082 => "0001100101001011",
4083 => "0001100101001100",4084 => "0001100101001100",
4085 => "0001100101001100",4086 => "0001100101001101",
4087 => "0001100101001101",4088 => "0001100101001101",
4089 => "0001100101001110",4090 => "0001100101001110",
4091 => "0001100101001110",4092 => "0001100101001111",
4093 => "0001100101001111",4094 => "0001100101001111",
4095 => "0001100101010000",4096 => "0011100110000101",
4097 => "0100000010100110",4098 => "0100100000011001",
4099 => "0100101111001110",4100 => "0101100000010111",
4101 => "0110000010110110",4102 => "0110100111010000",
4103 => "0111000001011000",4104 => "0000000000000000",
4105 => "0000000000000000",4106 => "0100000010100110",
4107 => "0100000011111000",4108 => "0100000101001011",
4109 => "0100000110011111",4110 => "0100000111110011",
4111 => "0100001001001001",4112 => "0100001010011111",
4113 => "0100001011110110",4114 => "0100001101001110",
4115 => "0100001110100111",4116 => "0100100000011001",
4117 => "0100100001110100",4118 => "0100100011001111",
4119 => "0100100000000011",4120 => "0100100110001001",
4121 => "0100100111101000",4122 => "0100101001000111",
4123 => "0100101010100111",4124 => "0100101100001001",
4125 => "0100101101101011",4126 => "0100101111001110",
4127 => "0101000001001010",4128 => "0101000010110000",
4129 => "0101000100010110",4130 => "0101000101111101",
4131 => "0101000111100110",4132 => "0101001001001111",
4133 => "0101001010111001",4134 => "0101001100100101",
4135 => "0101001110010001",4136 => "0101100000010111",
4137 => "0101100010000110",4138 => "0101100011110110",
4139 => "0101100101100111",4140 => "0101100111011001",
4141 => "0101101001001100",4142 => "0101101011000001",
4143 => "0101101100110110",4144 => "0101101110101101",
4145 => "0110000000111101",4146 => "0110000010110110",
4147 => "0110000100110001",4148 => "0110000110101101",
4149 => "0110001000101010",4150 => "0110000001000100",
4151 => "0110001100100111",4152 => "0110001110101000",
4153 => "0110100001000010",4154 => "0110100011000101",
4155 => "0110100000100001",4156 => "0110100111010000",
4157 => "0110101001010111",4158 => "0110101011100000",
4159 => "0110101101101010",4160 => "0111000000001101",
4161 => "0111000010011010",4162 => "0111000100101000",
4163 => "0111000000101100",4164 => "0111001001001001",
4165 => "0111001011011100",4166 => "0111000001011000",
4167 => "0111100000011101",4168 => "0111100000010010",
4169 => "0111100101001101",4170 => "0111100111100111",
4171 => "0000000000000000",4172 => "0000000000000000",
4173 => "0000000000000000",4174 => "0000000000000000",
4175 => "0000000000000000",4176 => "0000000000000000",
4177 => "0000000000000000",4178 => "0000000000000000",
4179 => "0000000000000000",4180 => "0000000000000000",
4181 => "0000000000000000",4182 => "0000000000000000",
4183 => "0000000000000000",4184 => "0000000000000000",
4185 => "0000000000000000",4186 => "0000000000000000",
4187 => "0000000000000000",4188 => "0000000000000000",
4189 => "0000000000000000",4190 => "0000000000000000",
4191 => "0000000000000000",4192 => "0000000000000000",
4193 => "0000000000000000",4194 => "0000000000000000",
4195 => "0000000000000000",4196 => "0100000010100110",
4197 => "0100000010101110",4198 => "0100000010110111",
4199 => "0100000010111111",4200 => "0100000011000111",
4201 => "0100000011001111",4202 => "0100000011010111",
4203 => "0100000011100000",4204 => "0100000011101000",
4205 => "0100000000011000",4206 => "0100000011111000",
4207 => "0100000100000000",4208 => "0100000100001001",
4209 => "0100000100010001",4210 => "0100000100011001",
4211 => "0100000000011101",4212 => "0100000100101010",
4213 => "0100000100110010",4214 => "0100000100111010",
4215 => "0100000101000011",4216 => "0100000101001011",
4217 => "0100000101010011",4218 => "0100000101011100",
4219 => "0100000101100100",4220 => "0100000101101101",
4221 => "0100000101110101",4222 => "0100000101111101",
4223 => "0100000000100111",4224 => "0100000110001110",
4225 => "0100000110010110",4226 => "0100000110011111",
4227 => "0100000110100111",4228 => "0100000110110000",
4229 => "0100000000101100",4230 => "0100000111000001",
4231 => "0100000111001001",4232 => "0100000111010010",
4233 => "0100000111011010",4234 => "0100000111100010",
4235 => "0100000111101011",4236 => "0100000111110011",
4237 => "0100000111111100",4238 => "0100001000000100",
4239 => "0100001000001101",4240 => "0100001000010110",
4241 => "0100001000011110",4242 => "0100001000100111",
4243 => "0100001000101111",4244 => "0100001000111000",
4245 => "0100001001000000",4246 => "0100001001001001",
4247 => "0100001001010001",4248 => "0100001001011010",
4249 => "0100001001100011",4250 => "0100001001101011",
4251 => "0100001001110100",4252 => "0100001001111101",
4253 => "0100001010000101",4254 => "0100001010001110",
4255 => "0100001010010110",4256 => "0100001010011111",
4257 => "0100000001000100",4258 => "0100001010110000",
4259 => "0100001010111001",4260 => "0100001011000010",
4261 => "0100001011001011",4262 => "0100001011010011",
4263 => "0100001011011100",4264 => "0100001011100101",
4265 => "0100000001001011",4266 => "0100001011110110",
4267 => "0100001011111111",4268 => "0100001100001000",
4269 => "0100001100010001",4270 => "0100001100011001",
4271 => "0100001100100010",4272 => "0100001100101011",
4273 => "0100000001010010",4274 => "0100001100111101",
4275 => "0100001101000101",4276 => "0100001101001110",
4277 => "0100001101010111",4278 => "0100001101100000",
4279 => "0100001101101001",4280 => "0100001101110010",
4281 => "0100001101111011",4282 => "0100000000001001",
4283 => "0100001110001100",4284 => "0100001110010101",
4285 => "0100001110011110",4286 => "0100001110100111",
4287 => "0100001110110000",4288 => "0100001110111001",
4289 => "0100001111000010",4290 => "0100001111001011",
4291 => "0100000001100010",4292 => "0100001111011101",
4293 => "0100001111100110",4294 => "0100100000000111",
4295 => "0100100000010000",4296 => "0100100000011001",
4297 => "0100100000100010",4298 => "0100100000101011",
4299 => "0100100000110100",4300 => "0100100000111101",
4301 => "0100100000000111",4302 => "0100100001001111",
4303 => "0100100001011000",4304 => "0100100001100010",
4305 => "0100100001101011",4306 => "0100100001110100",
4307 => "0100100001111101",4308 => "0100100010000110",
4309 => "0100100010001111",4310 => "0100100010011000",
4311 => "0100100010100001",4312 => "0100100010101011",
4313 => "0100100000010010",4314 => "0100100010111101",
4315 => "0100100011000110",4316 => "0100100011001111",
4317 => "0100100011011001",4318 => "0100100011100010",
4319 => "0100100011101011",4320 => "0100100011110100",
4321 => "0100100011111101",4322 => "0100100100000111",
4323 => "0100100100010000",4324 => "0100100100011001",
4325 => "0100100100100011",4326 => "0100100000000011",
4327 => "0100100100110101",4328 => "0100100100111110",
4329 => "0100100101001000",4330 => "0100100101010001",
4331 => "0100100101011010",4332 => "0100100101100100",
4333 => "0100100101101101",4334 => "0100100101110111",
4335 => "0100100110000000",4336 => "0100100110001001",
4337 => "0100100110010011",4338 => "0100100110011100",
4339 => "0100100110100110",4340 => "0100100110101111",
4341 => "0100100000101100",4342 => "0100100000101101",
4343 => "0100100111001011",4344 => "0100100111010101",
4345 => "0100100111011110",4346 => "0100100111101000",
4347 => "0100100111110001",4348 => "0100100111111011",
4349 => "0100101000000100",4350 => "0100101000001110",
4351 => "0100101000010111",4352 => "0100101000100001",
4353 => "0100101000101010",4354 => "0100101000110100",
4355 => "0100101000111110",4356 => "0100101001000111",
4357 => "0100101001010001",4358 => "0100101001011010",
4359 => "0100101001100100",4360 => "0100101001101101",
4361 => "0100101001110111",4362 => "0100101010000001",
4363 => "0100100001000001",4364 => "0100100001000010",
4365 => "0100100001000011",4366 => "0100101010100111",
4367 => "0100101010110001",4368 => "0100101010111011",
4369 => "0100101011000100",4370 => "0100101011001110",
4371 => "0100101011011000",4372 => "0100101011100010",
4373 => "0100101011101011",4374 => "0100101011110101",
4375 => "0100101011111111",4376 => "0100101100001001",
4377 => "0100101100010010",4378 => "0100101100011100",
4379 => "0100101100100110",4380 => "0100101100110000",
4381 => "0100101100111010",4382 => "0100101101000100",
4383 => "0100101101001101",4384 => "0100101101010111",
4385 => "0100101101100001",4386 => "0100101101101011",
4387 => "0100101101110101",4388 => "0100101101111111",
4389 => "0100101110001001",4390 => "0100101110010011",
4391 => "0100101110011100",4392 => "0100101110100110",
4393 => "0100101110110000",4394 => "0100101110111010",
4395 => "0100101111000100",4396 => "0100101111001110",
4397 => "0100101111011000",4398 => "0100101111100010",
4399 => "0101000000000100",4400 => "0101000000001110",
4401 => "0101000000011000",4402 => "0101000000100010",
4403 => "0101000000101100",4404 => "0101000000110110",
4405 => "0101000001000000",4406 => "0101000001001010",
4407 => "0101000001010101",4408 => "0101000001011111",
4409 => "0101000001101001",4410 => "0101000001110011",
4411 => "0101000001111101",4412 => "0101000010000111",
4413 => "0101000010010001",4414 => "0101000010011011",
4415 => "0101000010100110",4416 => "0101000010110000",
4417 => "0101000010111010",4418 => "0101000011000100",
4419 => "0101000011001110",4420 => "0101000011011000",
4421 => "0101000011100011",4422 => "0101000011101101",
4423 => "0101000011110111",4424 => "0101000100000001",
4425 => "0101000100001100",4426 => "0101000100010110",
4427 => "0101000100100000",4428 => "0101000100101011",
4429 => "0101000100110101",4430 => "0101000100111111",
4431 => "0101000101001001",4432 => "0101000000100010",
4433 => "0101000000100011",4434 => "0101000000100100",
4435 => "0101000101110011",4436 => "0101000101111101",
4437 => "0101000110001000",4438 => "0101000110010010",
4439 => "0101000110011100",4440 => "0101000110100111",
4441 => "0101000110110001",4442 => "0101000110111100",
4443 => "0101000111000110",4444 => "0101000111010001",
4445 => "0101000111011011",4446 => "0101000111100110",
4447 => "0101000111110000",4448 => "0101000111111011",
4449 => "0101001000000101",4450 => "0101001000010000",
4451 => "0101001000011010",4452 => "0101001000100101",
4453 => "0101001000101111",4454 => "0101000000111001",
4455 => "0101000000111010",4456 => "0101001001001111",
4457 => "0101001001011010",4458 => "0101001001100100",
4459 => "0101001001101111",4460 => "0101001001111001",
4461 => "0101001010000100",4462 => "0101001010001111",
4463 => "0101001010011001",4464 => "0101001010100100",
4465 => "0101001010101111",4466 => "0101001010111001",
4467 => "0101001011000100",4468 => "0101001011001111",
4469 => "0101000001001001",4470 => "0101000001001010",
4471 => "0101001011101111",4472 => "0101001011111010",
4473 => "0101001100000101",4474 => "0101001100001111",
4475 => "0101001100011010",4476 => "0101001100100101",
4477 => "0101001100110000",4478 => "0101001100111011",
4479 => "0101001101000101",4480 => "0101001101010000",
4481 => "0101001101011011",4482 => "0101000001010111",
4483 => "0101001101110001",4484 => "0101001101111100",
4485 => "0101001110000111",4486 => "0101001110010001",
4487 => "0101001110011100",4488 => "0101001110100111",
4489 => "0101001110110010",4490 => "0101001110111101",
4491 => "0101001111001000",4492 => "0101001111010011",
4493 => "0101000001100011",4494 => "0101100000000001",
4495 => "0101100000001100",4496 => "0101100000010111",
4497 => "0101100000100010",4498 => "0101100000101101",
4499 => "0101100000111000",4500 => "0101100001000011",
4501 => "0101100001001110",4502 => "0101100000001001",
4503 => "0101100001100101",4504 => "0101100001110000",
4505 => "0101100001111011",4506 => "0101100010000110",
4507 => "0101100010010001",4508 => "0101100010011100",
4509 => "0101100010100111",4510 => "0101100010110011",
4511 => "0101100000010011",4512 => "0101100011001001",
4513 => "0101100011010100",4514 => "0101100011011111",
4515 => "0101100011101011",4516 => "0101100011110110",
4517 => "0101100100000001",4518 => "0101100100001100",
4519 => "0101100000011100",4520 => "0101100100100011",
4521 => "0101100100101110",4522 => "0101100100111010",
4523 => "0101100101000101",4524 => "0101100101010000",
4525 => "0101100101011100",4526 => "0101100101100111",
4527 => "0101100000100101",4528 => "0101100101111110",
4529 => "0101100110001001",4530 => "0101100110010100",
4531 => "0101100110100000",4532 => "0101100110101011",
4533 => "0101100110110111",4534 => "0101100000101101",
4535 => "0101100111001110",4536 => "0101100111011001",
4537 => "0101100111100101",4538 => "0101100111110000",
4539 => "0101100111111100",4540 => "0101101000000111",
4541 => "0101101000010011",4542 => "0101101000011110",
4543 => "0101101000101010",4544 => "0101101000110101",
4545 => "0101101001000001",4546 => "0101101001001100",
4547 => "0101100000000110",4548 => "0101101001100100",
4549 => "0101101001101111",4550 => "0101101001111011",
4551 => "0101101010000110",4552 => "0101101010010010",
4553 => "0101100001000011",4554 => "0101101010101001",
4555 => "0101101010110101",4556 => "0101101011000001",
4557 => "0101101011001101",4558 => "0101101011011000",
4559 => "0101100001001010",4560 => "0101101011110000",
4561 => "0101101011111011",4562 => "0101101100000111",
4563 => "0101101100010011",4564 => "0101101100011111",
4565 => "0101101100101011",4566 => "0101101100110110",
4567 => "0101101101000010",4568 => "0101101101001110",
4569 => "0101101101011010",4570 => "0101100001010111",
4571 => "0101101101110010",4572 => "0101101101111110",
4573 => "0101101110001001",4574 => "0101101110010101",
4575 => "0101101110100001",4576 => "0101101110101101",
4577 => "0101101110111001",4578 => "0101101111000101",
4579 => "0101101111010001",4580 => "0101101111011101",
4581 => "0110000000000001",4582 => "0110000000001101",
4583 => "0110000000011001",4584 => "0110000000100101",
4585 => "0110000000110001",4586 => "0110000000111101",
4587 => "0110000001001001",4588 => "0110000001010101",
4589 => "0110000001100010",4590 => "0110000000001011",
4591 => "0110000001111010",4592 => "0110000010000110",
4593 => "0110000010010010",4594 => "0110000010011110",
4595 => "0110000000010001",4596 => "0110000010110110",
4597 => "0110000011000011",4598 => "0110000011001111",
4599 => "0110000011011011",4600 => "0110000011100111",
4601 => "0110000011110100",4602 => "0110000100000000",
4603 => "0110000100001100",4604 => "0110000000011100",
4605 => "0110000100100101",4606 => "0110000100110001",
4607 => "0110000100111101",4608 => "0110000000100001",
4609 => "0110000101010110",4610 => "0110000101100010",
4611 => "0110000101101111",4612 => "0110000101111011",
4613 => "0110000110000111",4614 => "0110000110010100",
4615 => "0110000110100000",4616 => "0110000110101101",
4617 => "0110000110111001",4618 => "0110000111000101",
4619 => "0110000111010010",4620 => "0110000111011110",
4621 => "0110000111101011",4622 => "0110000111110111",
4623 => "0110001000000100",4624 => "0110001000010000",
4625 => "0110001000011101",4626 => "0110001000101010",
4627 => "0110001000110110",4628 => "0110001001000011",
4629 => "0110001001001111",4630 => "0110001001011100",
4631 => "0110001001101000",4632 => "0110001001110101",
4633 => "0110001010000010",4634 => "0110001010001110",
4635 => "0110001010011011",4636 => "0110000001000100",
4637 => "0110001010110100",4638 => "0110001011000001",
4639 => "0110001011001110",4640 => "0110000001001001",
4641 => "0110001011100111",4642 => "0110001011110100",
4643 => "0110001100000001",4644 => "0110001100001110",
4645 => "0110001100011010",4646 => "0110001100100111",
4647 => "0110000001010010",4648 => "0110001101000001",
4649 => "0110001101001110",4650 => "0110001101011010",
4651 => "0110001101100111",4652 => "0110001101110100",
4653 => "0110001110000001",4654 => "0110000001011011",
4655 => "0110001110011011",4656 => "0110001110101000",
4657 => "0110001110110101",4658 => "0110001111000010",
4659 => "0110001111001111",4660 => "0110001111011100",
4661 => "0110100000000001",4662 => "0110100000001110",
4663 => "0110100000011011",4664 => "0110100000000100",
4665 => "0110100000110101",4666 => "0110100001000010",
4667 => "0110100001001111",4668 => "0110100001011100",
4669 => "0110100001101001",4670 => "0110100001110110",
4671 => "0110100010000011",4672 => "0110100010010000",
4673 => "0110100010011110",4674 => "0110100010101011",
4675 => "0110100010111000",4676 => "0110100011000101",
4677 => "0110100000010101",4678 => "0110100011100000",
4679 => "0110100011101101",4680 => "0110100000011001",
4681 => "0110100100000111",4682 => "0110100100010101",
4683 => "0110100000011101",4684 => "0110100100101111",
4685 => "0110100100111100",4686 => "0110100000100001",
4687 => "0110100101010111",4688 => "0110100101100100",
4689 => "0110100000100101",4690 => "0110100101111111",
4691 => "0110100110001101",4692 => "0110100000101001",
4693 => "0110100110100111",4694 => "0110100110110101",
4695 => "0110100000101101",4696 => "0110100111010000",
4697 => "0110100111011101",4698 => "0110100111101011",
4699 => "0110100111111000",4700 => "0110101000000110",
4701 => "0110101000010011",4702 => "0110101000100001",
4703 => "0110101000101110",4704 => "0110101000111100",
4705 => "0110101001001001",4706 => "0110101001010111",
4707 => "0110101001100101",4708 => "0110101001110010",
4709 => "0110100001000000",4710 => "0110101010001110",
4711 => "0110101010011011",4712 => "0110101010101001",
4713 => "0110101010110111",4714 => "0110101011000100",
4715 => "0110101011010010",4716 => "0110101011100000",
4717 => "0110101011101101",4718 => "0110101011111011",
4719 => "0110101100001001",4720 => "0110101100010111",
4721 => "0110101100100101",4722 => "0110101100110010",
4723 => "0110101101000000",4724 => "0110101101001110",
4725 => "0110100001010110",4726 => "0110101101101010",
4727 => "0110101101111000",4728 => "0110101110000110",
4729 => "0110101110010011",4730 => "0110101110100001",
4731 => "0110101110101111",4732 => "0110101110111101",
4733 => "0110101111001011",4734 => "0110101111011001",
4735 => "0110101111100111",4736 => "0111000000001101",
4737 => "0111000000011011",4738 => "0111000000101001",
4739 => "0111000000110111",4740 => "0111000001000101",
4741 => "0111000001010011",4742 => "0111000001100010",
4743 => "0111000001110000",4744 => "0111000001111110",
4745 => "0111000000001110",4746 => "0111000010011010",
4747 => "0111000010101000",4748 => "0111000010110110",
4749 => "0111000011000101",4750 => "0111000011010011",
4751 => "0111000011100001",4752 => "0111000011101111",
4753 => "0111000011111101",4754 => "0111000100001100",
4755 => "0111000100011010",4756 => "0111000100101000",
4757 => "0111000100110111",4758 => "0111000101000101",
4759 => "0111000101010011",4760 => "0111000101100010",
4761 => "0111000101110000",4762 => "0111000101111110",
4763 => "0111000110001101",4764 => "0111000110011011",
4765 => "0111000110101010",4766 => "0111000000101100",
4767 => "0111000111000110",4768 => "0111000111010101",
4769 => "0111000111100011",4770 => "0111000111110010",
4771 => "0111001000000000",4772 => "0111001000001111",
4773 => "0111001000011101",4774 => "0111001000101100",
4775 => "0111001000111011",4776 => "0111001001001001",
4777 => "0111000000000110",4778 => "0111001001100110",
4779 => "0111001001110101",4780 => "0111001010000100",
4781 => "0111001010010010",4782 => "0111001010100001",
4783 => "0111001010110000",4784 => "0111001010111110",
4785 => "0111001011001101",4786 => "0111001011011100",
4787 => "0111001011101010",4788 => "0111001011111001",
4789 => "0111001100001000",4790 => "0111001100010111",
4791 => "0111001100100110",4792 => "0111000001010010",
4793 => "0111001101000011",4794 => "0111000001010101",
4795 => "0111001101100001",4796 => "0111000001011000",
4797 => "0111001101111111",4798 => "0111000001011011",
4799 => "0111001110011100",4800 => "0111001110101011",
4801 => "0111001110111010",4802 => "0111001111001001",
4803 => "0111001111011000",4804 => "0111001111100111",
4805 => "0111100000001110",4806 => "0111100000011101",
4807 => "0111100000101100",4808 => "0111100000111011",
4809 => "0111100001001010",4810 => "0111100000001001",
4811 => "0111100001101001",4812 => "0111100000001100",
4813 => "0111100010000111",4814 => "0111100000001111",
4815 => "0111100010100101",4816 => "0111100000010010",
4817 => "0111100011000100",4818 => "0111100011010011",
4819 => "0111100011100010",4820 => "0111100011110001",
4821 => "0111100100000000",4822 => "0111100100010000",
4823 => "0111100100011111",4824 => "0111100100101110",
4825 => "0111100100111110",4826 => "0111100101001101",
4827 => "0111100101011100",4828 => "0111100101101100",
4829 => "0111100101111011",4830 => "0111100110001010",
4831 => "0111100000101001",4832 => "0111100110101001",
4833 => "0111100110111001",4834 => "0111100111001000",
4835 => "0111100111011000",4836 => "0111100111100111",
4837 => "0000000000000000",4838 => "0000000000000000",
4839 => "0000000000000000",4840 => "0000000000000000",
4841 => "0000000000000000",4842 => "0000000000000000",
4843 => "0000000000000000",4844 => "0000000000000000",
4845 => "0000000000000000",4846 => "0000000000000000",
4847 => "0000000000000000",4848 => "0000000000000000",
4849 => "0000000000000000",4850 => "0000000000000000",
4851 => "0000000000000000",4852 => "0000000000000000",
4853 => "0000000000000000",4854 => "0000000000000000",
4855 => "0000000000000000",4856 => "0000000000000000",
4857 => "0000000000000000",4858 => "0000000000000000",
4859 => "0000000000000000",4860 => "0000000000000000",
4861 => "0000000000000000",4862 => "0000000000000000",
4863 => "0000000000000000",4864 => "0000000000000000",
4865 => "0000000000000000",4866 => "0000000000000000",
4867 => "0000000000000000",4868 => "0000000000000000",
4869 => "0000000000000000",4870 => "0000000000000000",
4871 => "0000000000000000",4872 => "0000000000000000",
4873 => "0000000000000000",4874 => "0000000000000000",
4875 => "0000000000000000",4876 => "0000000000000000",
4877 => "0000000000000000",4878 => "0000000000000000",
4879 => "0000000000000000",4880 => "0000000000000000",
4881 => "0000000000000000",4882 => "0000000000000000",
4883 => "0000000000000000",4884 => "0000000000000000",
4885 => "0000000000000000",4886 => "0000000000000000",
4887 => "0000000000000000",4888 => "0000000000000000",
4889 => "0000000000000000",4890 => "0000000000000000",
4891 => "0000000000000000",4892 => "0000000000000000",
4893 => "0000000000000000",4894 => "0000000000000000",
4895 => "0000000000000000",4896 => "0000000000000000",
4897 => "0000000000000000",4898 => "0000000000000000",
4899 => "0000000000000000",4900 => "0000000000000000",
4901 => "0000000000000000",4902 => "0000000000000000",
4903 => "0000000000000000",4904 => "0000000000000000",
4905 => "0000000000000000",4906 => "0000000000000000",
4907 => "0000000000000000",4908 => "0000000000000000",
4909 => "0000000000000000",4910 => "0000000000000000",
4911 => "0000000000000000",4912 => "0000000000000000",
4913 => "0000000000000000",4914 => "0000000000000000",
4915 => "0000000000000000",4916 => "0000000000000000",
4917 => "0000000000000000",4918 => "0000000000000000",
4919 => "0000000000000000",4920 => "0000000000000000",
4921 => "0000000000000000",4922 => "0000000000000000",
4923 => "0000000000000000",4924 => "0000000000000000",
4925 => "0000000000000000",4926 => "0000000000000000",
4927 => "0000000000000000",4928 => "0000000000000000",
4929 => "0000000000000000",4930 => "0000000000000000",
4931 => "0000000000000000",4932 => "0000000000000000",
4933 => "0000000000000000",4934 => "0000000000000000",
4935 => "0000000000000000",4936 => "0000000000000000",
4937 => "0000000000000000",4938 => "0000000000000000",
4939 => "0000000000000000",4940 => "0000000000000000",
4941 => "0000000000000000",4942 => "0000000000000000",
4943 => "0000000000000000",4944 => "0000000000000000",
4945 => "0000000000000000",4946 => "0000000000000000",
4947 => "0000000000000000",4948 => "0000000000000000",
4949 => "0000000000000000",4950 => "0000000000000000",
4951 => "0000000000000000",4952 => "0000000000000000",
4953 => "0000000000000000",4954 => "0000000000000000",
4955 => "0000000000000000",4956 => "0000000000000000",
4957 => "0000000000000000",4958 => "0000000000000000",
4959 => "0000000000000000",4960 => "0000000000000000",
4961 => "0000000000000000",4962 => "0000000000000000",
4963 => "0000000000000000",4964 => "0000000000000000",
4965 => "0000000000000000",4966 => "0000000000000000",
4967 => "0000000000000000",4968 => "0000000000000000",
4969 => "0000000000000000",4970 => "0000000000000000",
4971 => "0000000000000000",4972 => "0000000000000000",
4973 => "0000000000000000",4974 => "0000000000000000",
4975 => "0000000000000000",4976 => "0000000000000000",
4977 => "0000000000000000",4978 => "0000000000000000",
4979 => "0000000000000000",4980 => "0000000000000000",
4981 => "0000000000000000",4982 => "0000000000000000",
4983 => "0000000000000000",4984 => "0000000000000000",
4985 => "0000000000000000",4986 => "0000000000000000",
4987 => "0000000000000000",4988 => "0000000000000000",
4989 => "0000000000000000",4990 => "0000000000000000",
4991 => "0000000000000000",4992 => "0000000000000000",
4993 => "0000000000000000",4994 => "0000000000000000",
4995 => "0000000000000000",4996 => "0000000000000000",
4997 => "0000000000000000",4998 => "0000000000000000",
4999 => "0000000000000000",5000 => "0000000000000000",
5001 => "0000000000000000",5002 => "0000000000000000",
5003 => "0000000000000000",5004 => "0000000000000000",
5005 => "0000000000000000",5006 => "0000000000000000",
5007 => "0000000000000000",5008 => "0000000000000000",
5009 => "0000000000000000",5010 => "0000000000000000",
5011 => "0000000000000000",5012 => "0000000000000000",
5013 => "0000000000000000",5014 => "0000000000000000",
5015 => "0000000000000000",5016 => "0000000000000000",
5017 => "0000000000000000",5018 => "0000000000000000",
5019 => "0000000000000000",5020 => "0000000000000000",
5021 => "0000000000000000",5022 => "0000000000000000",
5023 => "0000000000000000",5024 => "0000000000000000",
5025 => "0000000000000000",5026 => "0000000000000000",
5027 => "0000000000000000",5028 => "0000000000000000",
5029 => "0000000000000000",5030 => "0000000000000000",
5031 => "0000000000000000",5032 => "0000000000000000",
5033 => "0000000000000000",5034 => "0000000000000000",
5035 => "0000000000000000",5036 => "0000000000000000",
5037 => "0000000000000000",5038 => "0000000000000000",
5039 => "0000000000000000",5040 => "0000000000000000",
5041 => "0000000000000000",5042 => "0000000000000000",
5043 => "0000000000000000",5044 => "0000000000000000",
5045 => "0000000000000000",5046 => "0000000000000000",
5047 => "0000000000000000",5048 => "0000000000000000",
5049 => "0000000000000000",5050 => "0000000000000000",
5051 => "0000000000000000",5052 => "0000000000000000",
5053 => "0000000000000000",5054 => "0000000000000000",
5055 => "0000000000000000",5056 => "0000000000000000",
5057 => "0000000000000000",5058 => "0000000000000000",
5059 => "0000000000000000",5060 => "0000000000000000",
5061 => "0000000000000000",5062 => "0000000000000000",
5063 => "0000000000000000",5064 => "0000000000000000",
5065 => "0000000000000000",5066 => "0000000000000000",
5067 => "0000000000000000",5068 => "0000000000000000",
5069 => "0000000000000000",5070 => "0000000000000000",
5071 => "0000000000000000",5072 => "0000000000000000",
5073 => "0000000000000000",5074 => "0000000000000000",
5075 => "0000000000000000",5076 => "0000000000000000",
5077 => "0000000000000000",5078 => "0000000000000000",
5079 => "0000000000000000",5080 => "0000000000000000",
5081 => "0000000000000000",5082 => "0000000000000000",
5083 => "0000000000000000",5084 => "0000000000000000",
5085 => "0000000000000000",5086 => "0000000000000000",
5087 => "0000000000000000",5088 => "0000000000000000",
5089 => "0000000000000000",5090 => "0000000000000000",
5091 => "0000000000000000",5092 => "0000000000000000",
5093 => "0000000000000000",5094 => "0000000000000000",
5095 => "0000000000000000",5096 => "0100000010100110",
5097 => "0100000010100111",5098 => "0100000010101000",
5099 => "0100000010101001",5100 => "0100000010101001",
5101 => "0100000000010001",5102 => "0100000010101011",
5103 => "0100000010101100",5104 => "0100000010101101",
5105 => "0100000010101110",5106 => "0100000010101110",
5107 => "0100000010101111",5108 => "0100000010110000",
5109 => "0100000010110001",5110 => "0100000010110010",
5111 => "0100000010110010",5112 => "0100000010110011",
5113 => "0100000000010010",5114 => "0100000010110101",
5115 => "0100000010110110",5116 => "0100000010110111",
5117 => "0100000010110111",5118 => "0100000010111000",
5119 => "0100000010111001",5120 => "0100000010111010",
5121 => "0100000010111011",5122 => "0100000010111011",
5123 => "0100000010111100",5124 => "0100000010111101",
5125 => "0100000000010011",5126 => "0100000010111111",
5127 => "0100000011000000",5128 => "0100000011000000",
5129 => "0100000011000001",5130 => "0100000011000010",
5131 => "0100000011000011",5132 => "0100000011000100",
5133 => "0100000011000100",5134 => "0100000011000101",
5135 => "0100000011000110",5136 => "0100000011000111",
5137 => "0100000000000010",5138 => "0100000011001001",
5139 => "0100000011001001",5140 => "0100000011001010",
5141 => "0100000011001011",5142 => "0100000011001100",
5143 => "0100000011001101",5144 => "0100000011001101",
5145 => "0100000011001110",5146 => "0100000011001111",
5147 => "0100000011010000",5148 => "0100000011010001",
5149 => "0100000000010101",5150 => "0100000000010101",
5151 => "0100000011010011",5152 => "0100000011010100",
5153 => "0100000011010101",5154 => "0100000011010110",
5155 => "0100000011010110",5156 => "0100000011010111",
5157 => "0100000011011000",5158 => "0100000011011001",
5159 => "0100000011011010",5160 => "0100000011011011",
5161 => "0100000011011011",5162 => "0100000000010110",
5163 => "0100000011011101",5164 => "0100000011011110",
5165 => "0100000011011111",5166 => "0100000011100000",
5167 => "0100000011100000",5168 => "0100000011100001",
5169 => "0100000011100010",5170 => "0100000011100011",
5171 => "0100000011100100",5172 => "0100000011100100",
5173 => "0100000011100101",5174 => "0100000000010111",
5175 => "0100000011100111",5176 => "0100000011101000",
5177 => "0100000011101001",5178 => "0100000011101001",
5179 => "0100000011101010",5180 => "0100000011101011",
5181 => "0100000011101100",5182 => "0100000011101101",
5183 => "0100000011101110",5184 => "0100000011101110",
5185 => "0100000011101111",5186 => "0100000000011000",
5187 => "0100000011110001",5188 => "0100000011110010",
5189 => "0100000011110010",5190 => "0100000011110011",
5191 => "0100000011110100",5192 => "0100000011110101",
5193 => "0100000011110110",5194 => "0100000011110111",
5195 => "0100000011110111",5196 => "0100000011111000",
5197 => "0100000011111001",5198 => "0100000000011001",
5199 => "0100000011111011",5200 => "0100000011111100",
5201 => "0100000011111100",5202 => "0100000011111101",
5203 => "0100000011111110",5204 => "0100000011111111",
5205 => "0100000100000000",5206 => "0100000100000000",
5207 => "0100000100000001",5208 => "0100000100000010",
5209 => "0100000100000011",5210 => "0100000000011010",
5211 => "0100000100000101",5212 => "0100000100000101",
5213 => "0100000100000110",5214 => "0100000100000111",
5215 => "0100000100001000",5216 => "0100000100001001",
5217 => "0100000100001010",5218 => "0100000100001010",
5219 => "0100000100001011",5220 => "0100000100001100",
5221 => "0100000100001101",5222 => "0100000000011011",
5223 => "0100000100001111",5224 => "0100000100001111",
5225 => "0100000100010000",5226 => "0100000100010001",
5227 => "0100000100010010",5228 => "0100000100010011",
5229 => "0100000100010100",5230 => "0100000100010100",
5231 => "0100000100010101",5232 => "0100000100010110",
5233 => "0100000100010111",5234 => "0100000000011100",
5235 => "0100000000011100",5236 => "0100000100011001",
5237 => "0100000100011010",5238 => "0100000100011011",
5239 => "0100000100011100",5240 => "0100000100011101",
5241 => "0100000100011101",5242 => "0100000100011110",
5243 => "0100000100011111",5244 => "0100000100100000",
5245 => "0100000100100001",5246 => "0100000000011101",
5247 => "0100000000011101",5248 => "0100000100100011",
5249 => "0100000100100100",5250 => "0100000100100101",
5251 => "0100000100100110",5252 => "0100000100100111",
5253 => "0100000100100111",5254 => "0100000100101000",
5255 => "0100000100101001",5256 => "0100000100101010",
5257 => "0100000100101011",5258 => "0100000000000011",
5259 => "0100000000000011",5260 => "0100000100101101",
5261 => "0100000100101110",5262 => "0100000100101111",
5263 => "0100000100110000",5264 => "0100000100110001",
5265 => "0100000100110001",5266 => "0100000100110010",
5267 => "0100000100110011",5268 => "0100000100110100",
5269 => "0100000100110101",5270 => "0100000000011111",
5271 => "0100000000011111",5272 => "0100000100110111",
5273 => "0100000100111000",5274 => "0100000100111001",
5275 => "0100000100111010",5276 => "0100000100111010",
5277 => "0100000100111011",5278 => "0100000100111100",
5279 => "0100000100111101",5280 => "0100000100111110",
5281 => "0100000100111111",5282 => "0100000100111111",
5283 => "0100000000100000",5284 => "0100000101000001",
5285 => "0100000101000010",5286 => "0100000101000011",
5287 => "0100000101000100",5288 => "0100000101000100",
5289 => "0100000101000101",5290 => "0100000101000110",
5291 => "0100000101000111",5292 => "0100000101001000",
5293 => "0100000101001001",5294 => "0100000101001001",
5295 => "0100000000100001",5296 => "0100000101001011",
5297 => "0100000101001100",5298 => "0100000101001101",
5299 => "0100000101001110",5300 => "0100000101001110",
5301 => "0100000101001111",5302 => "0100000101010000",
5303 => "0100000101010001",5304 => "0100000101010010",
5305 => "0100000101010011",5306 => "0100000101010011",
5307 => "0100000000100010",5308 => "0100000101010101",
5309 => "0100000101010110",5310 => "0100000101010111",
5311 => "0100000101011000",5312 => "0100000101011000",
5313 => "0100000101011001",5314 => "0100000101011010",
5315 => "0100000101011011",5316 => "0100000101011100",
5317 => "0100000101011101",5318 => "0100000101011101",
5319 => "0100000000100011",5320 => "0100000101011111",
5321 => "0100000101100000",5322 => "0100000101100001",
5323 => "0100000101100010",5324 => "0100000101100010",
5325 => "0100000101100011",5326 => "0100000101100100",
5327 => "0100000101100101",5328 => "0100000101100110",
5329 => "0100000101100111",5330 => "0100000000100100",
5331 => "0100000000100100",5332 => "0100000101101001",
5333 => "0100000101101010",5334 => "0100000101101011",
5335 => "0100000101101100",5336 => "0100000101101101",
5337 => "0100000101101101",5338 => "0100000101101110",
5339 => "0100000101101111",5340 => "0100000101110000",
5341 => "0100000101110001",5342 => "0100000000100101",
5343 => "0100000000100101",5344 => "0100000101110011",
5345 => "0100000101110100",5346 => "0100000101110101",
5347 => "0100000101110110",5348 => "0100000101110111",
5349 => "0100000101110111",5350 => "0100000101111000",
5351 => "0100000101111001",5352 => "0100000101111010",
5353 => "0100000101111011",5354 => "0100000000100110",
5355 => "0100000000100110",5356 => "0100000101111101",
5357 => "0100000101111110",5358 => "0100000101111111",
5359 => "0100000110000000",5360 => "0100000110000001",
5361 => "0100000110000001",5362 => "0100000110000010",
5363 => "0100000110000011",5364 => "0100000110000100",
5365 => "0100000110000101",5366 => "0100000000100111",
5367 => "0100000000100111",5368 => "0100000110000111",
5369 => "0100000110001000",5370 => "0100000110001001",
5371 => "0100000110001010",5372 => "0100000110001011",
5373 => "0100000110001100",5374 => "0100000110001100",
5375 => "0100000110001101",5376 => "0100000110001110",
5377 => "0100000110001111",5378 => "0100000000000100",
5379 => "0100000110010001",5380 => "0100000110010001",
5381 => "0100000110010010",5382 => "0100000110010011",
5383 => "0100000110010100",5384 => "0100000110010101",
5385 => "0100000110010110",5386 => "0100000110010110",
5387 => "0100000110010111",5388 => "0100000110011000",
5389 => "0100000110011001",5390 => "0100000000101001",
5391 => "0100000110011011",5392 => "0100000110011100",
5393 => "0100000110011100",5394 => "0100000110011101",
5395 => "0100000110011110",5396 => "0100000110011111",
5397 => "0100000110100000",5398 => "0100000110100001",
5399 => "0100000110100001",5400 => "0100000110100010",
5401 => "0100000110100011",5402 => "0100000000101010",
5403 => "0100000110100101",5404 => "0100000110100110",
5405 => "0100000110100110",5406 => "0100000110100111",
5407 => "0100000110101000",5408 => "0100000110101001",
5409 => "0100000110101010",5410 => "0100000110101011",
5411 => "0100000110101011",5412 => "0100000110101100",
5413 => "0100000110101101",5414 => "0100000000101011",
5415 => "0100000110101111",5416 => "0100000110110000",
5417 => "0100000110110001",5418 => "0100000110110001",
5419 => "0100000110110010",5420 => "0100000110110011",
5421 => "0100000110110100",5422 => "0100000110110101",
5423 => "0100000110110110",5424 => "0100000110110110",
5425 => "0100000110110111",5426 => "0100000000101100",
5427 => "0100000110111001",5428 => "0100000110111010",
5429 => "0100000110111011",5430 => "0100000110111100",
5431 => "0100000110111100",5432 => "0100000110111101",
5433 => "0100000110111110",5434 => "0100000110111111",
5435 => "0100000111000000",5436 => "0100000111000001",
5437 => "0100000111000001",5438 => "0100000000101101",
5439 => "0100000111000011",5440 => "0100000111000100",
5441 => "0100000111000101",5442 => "0100000111000110",
5443 => "0100000111000111",5444 => "0100000111000111",
5445 => "0100000111001000",5446 => "0100000111001001",
5447 => "0100000111001010",5448 => "0100000111001011",
5449 => "0100000000101110",5450 => "0100000000101110",
5451 => "0100000111001101",5452 => "0100000111001110",
5453 => "0100000111001111",5454 => "0100000111010000",
5455 => "0100000111010001",5456 => "0100000111010010",
5457 => "0100000111010010",5458 => "0100000111010011",
5459 => "0100000111010100",5460 => "0100000111010101",
5461 => "0100000000101111",5462 => "0100000111010111",
5463 => "0100000111010111",5464 => "0100000111011000",
5465 => "0100000111011001",5466 => "0100000111011010",
5467 => "0100000111011011",5468 => "0100000111011100",
5469 => "0100000111011101",5470 => "0100000111011101",
5471 => "0100000111011110",5472 => "0100000111011111",
5473 => "0100000000110000",5474 => "0100000111100001",
5475 => "0100000111100010",5476 => "0100000111100010",
5477 => "0100000111100011",5478 => "0100000111100100",
5479 => "0100000111100101",5480 => "0100000111100110",
5481 => "0100000111100111",5482 => "0100000111101000",
5483 => "0100000111101000",5484 => "0100000111101001",
5485 => "0100000000110001",5486 => "0100000111101011",
5487 => "0100000111101100",5488 => "0100000111101101",
5489 => "0100000111101101",5490 => "0100000111101110",
5491 => "0100000111101111",5492 => "0100000111110000",
5493 => "0100000111110001",5494 => "0100000111110010",
5495 => "0100000111110011",5496 => "0100000111110011",
5497 => "0100000000000101",5498 => "0100000111110101",
5499 => "0100000111110110",5500 => "0100000111110111",
5501 => "0100000111111000",5502 => "0100000111111001",
5503 => "0100000111111001",5504 => "0100000111111010",
5505 => "0100000111111011",5506 => "0100000111111100",
5507 => "0100000111111101",5508 => "0100000000110011",
5509 => "0100000000110011",5510 => "0100000111111111",
5511 => "0100001000000000",5512 => "0100001000000001",
5513 => "0100001000000010",5514 => "0100001000000011",
5515 => "0100001000000100",5516 => "0100001000000100",
5517 => "0100001000000101",5518 => "0100001000000110",
5519 => "0100001000000111",5520 => "0100000000110100",
5521 => "0100001000001001",5522 => "0100001000001010",
5523 => "0100001000001010",5524 => "0100001000001011",
5525 => "0100001000001100",5526 => "0100001000001101",
5527 => "0100001000001110",5528 => "0100001000001111",
5529 => "0100001000010000",5530 => "0100001000010000",
5531 => "0100001000010001",5532 => "0100000000110101",
5533 => "0100001000010011",5534 => "0100001000010100",
5535 => "0100001000010101",5536 => "0100001000010110",
5537 => "0100001000010110",5538 => "0100001000010111",
5539 => "0100001000011000",5540 => "0100001000011001",
5541 => "0100001000011010",5542 => "0100001000011011",
5543 => "0100001000011011",5544 => "0100000000110110",
5545 => "0100001000011101",5546 => "0100001000011110",
5547 => "0100001000011111",5548 => "0100001000100000",
5549 => "0100001000100001",5550 => "0100001000100001",
5551 => "0100001000100010",5552 => "0100001000100011",
5553 => "0100001000100100",5554 => "0100001000100101",
5555 => "0100000000110111",5556 => "0100001000100111",
5557 => "0100001000100111",5558 => "0100001000101000",
5559 => "0100001000101001",5560 => "0100001000101010",
5561 => "0100001000101011",5562 => "0100001000101100",
5563 => "0100001000101101",5564 => "0100001000101101",
5565 => "0100001000101110",5566 => "0100001000101111",
5567 => "0100000000111000",5568 => "0100001000110001",
5569 => "0100001000110010",5570 => "0100001000110011",
5571 => "0100001000110011",5572 => "0100001000110100",
5573 => "0100001000110101",5574 => "0100001000110110",
5575 => "0100001000110111",5576 => "0100001000111000",
5577 => "0100001000111001",5578 => "0100001000111001",
5579 => "0100000000111001",5580 => "0100001000111011",
5581 => "0100001000111100",5582 => "0100001000111101",
5583 => "0100001000111110",5584 => "0100001000111111",
5585 => "0100001000111111",5586 => "0100001001000000",
5587 => "0100001001000001",5588 => "0100001001000010",
5589 => "0100001001000011",5590 => "0100000000111010",
5591 => "0100001001000101",5592 => "0100001001000101",
5593 => "0100001001000110",5594 => "0100001001000111",
5595 => "0100001001001000",5596 => "0100001001001001",
5597 => "0100001001001010",5598 => "0100001001001011",
5599 => "0100001001001011",5600 => "0100001001001100",
5601 => "0100001001001101",5602 => "0100000000111011",
5603 => "0100001001001111",5604 => "0100001001010000",
5605 => "0100001001010001",5606 => "0100001001010001",
5607 => "0100001001010010",5608 => "0100001001010011",
5609 => "0100001001010100",5610 => "0100001001010101",
5611 => "0100001001010110",5612 => "0100001001010111",
5613 => "0100001001010111",5614 => "0100000000000110",
5615 => "0100001001011001",5616 => "0100001001011010",
5617 => "0100001001011011",5618 => "0100001001011100",
5619 => "0100001001011101",5620 => "0100001001011101",
5621 => "0100001001011110",5622 => "0100001001011111",
5623 => "0100001001100000",5624 => "0100001001100001",
5625 => "0100000000111101",5626 => "0100001001100011",
5627 => "0100001001100100",5628 => "0100001001100100",
5629 => "0100001001100101",5630 => "0100001001100110",
5631 => "0100001001100111",5632 => "0100001001101000",
5633 => "0100001001101001",5634 => "0100001001101010",
5635 => "0100001001101010",5636 => "0100001001101011",
5637 => "0100000000111110",5638 => "0100001001101101",
5639 => "0100001001101110",5640 => "0100001001101111",
5641 => "0100001001110000",5642 => "0100001001110000",
5643 => "0100001001110001",5644 => "0100001001110010",
5645 => "0100001001110011",5646 => "0100001001110100",
5647 => "0100001001110101",5648 => "0100000000111111",
5649 => "0100000000111111",5650 => "0100001001110111",
5651 => "0100001001111000",5652 => "0100001001111001",
5653 => "0100001001111010",5654 => "0100001001111011",
5655 => "0100001001111100",5656 => "0100001001111101",
5657 => "0100001001111101",5658 => "0100001001111110",
5659 => "0100001001111111",5660 => "0100000001000000",
5661 => "0100001010000001",5662 => "0100001010000010",
5663 => "0100001010000011",5664 => "0100001010000011",
5665 => "0100001010000100",5666 => "0100001010000101",
5667 => "0100001010000110",5668 => "0100001010000111",
5669 => "0100001010001000",5670 => "0100001010001001",
5671 => "0100001010001001",5672 => "0100000001000001",
5673 => "0100001010001011",5674 => "0100001010001100",
5675 => "0100001010001101",5676 => "0100001010001110",
5677 => "0100001010001111",5678 => "0100001010010000",
5679 => "0100001010010000",5680 => "0100001010010001",
5681 => "0100001010010010",5682 => "0100001010010011",
5683 => "0100000001000010",5684 => "0100001010010101",
5685 => "0100001010010110",5686 => "0100001010010110",
5687 => "0100001010010111",5688 => "0100001010011000",
5689 => "0100001010011001",5690 => "0100001010011010",
5691 => "0100001010011011",5692 => "0100001010011100",
5693 => "0100001010011101",5694 => "0100001010011101",
5695 => "0100000001000011",5696 => "0100001010011111",
5697 => "0100001010100000",5698 => "0100001010100001",
5699 => "0100001010100010",5700 => "0100001010100011",
5701 => "0100001010100011",5702 => "0100001010100100",
5703 => "0100001010100101",5704 => "0100001010100110",
5705 => "0100001010100111",5706 => "0100000001000100",
5707 => "0100001010101001",5708 => "0100001010101010",
5709 => "0100001010101010",5710 => "0100001010101011",
5711 => "0100001010101100",5712 => "0100001010101101",
5713 => "0100001010101110",5714 => "0100001010101111",
5715 => "0100001010110000",5716 => "0100001010110000",
5717 => "0100001010110001",5718 => "0100000001000101",
5719 => "0100001010110011",5720 => "0100001010110100",
5721 => "0100001010110101",5722 => "0100001010110110",
5723 => "0100001010110111",5724 => "0100001010110111",
5725 => "0100001010111000",5726 => "0100001010111001",
5727 => "0100001010111010",5728 => "0100001010111011",
5729 => "0100000000000111",5730 => "0100001010111101",
5731 => "0100001010111110",5732 => "0100001010111110",
5733 => "0100001010111111",5734 => "0100001011000000",
5735 => "0100001011000001",5736 => "0100001011000010",
5737 => "0100001011000011",5738 => "0100001011000100",
5739 => "0100001011000101",5740 => "0100001011000101",
5741 => "0100000001000111",5742 => "0100001011000111",
5743 => "0100001011001000",5744 => "0100001011001001",
5745 => "0100001011001010",5746 => "0100001011001011",
5747 => "0100001011001011",5748 => "0100001011001100",
5749 => "0100001011001101",5750 => "0100001011001110",
5751 => "0100001011001111",5752 => "0100000001001000",
5753 => "0100001011010001",5754 => "0100001011010010",
5755 => "0100001011010010",5756 => "0100001011010011",
5757 => "0100001011010100",5758 => "0100001011010101",
5759 => "0100001011010110",5760 => "0100001011010111",
5761 => "0100001011011000",5762 => "0100001011011001",
5763 => "0100001011011001",5764 => "0100000001001001",
5765 => "0100001011011011",5766 => "0100001011011100",
5767 => "0100001011011101",5768 => "0100001011011110",
5769 => "0100001011011111",5770 => "0100001011100000",
5771 => "0100001011100000",5772 => "0100001011100001",
5773 => "0100001011100010",5774 => "0100001011100011",
5775 => "0100000001001010",5776 => "0100001011100101",
5777 => "0100001011100110",5778 => "0100001011100111",
5779 => "0100001011100111",5780 => "0100001011101000",
5781 => "0100001011101001",5782 => "0100001011101010",
5783 => "0100001011101011",5784 => "0100001011101100",
5785 => "0100001011101101",5786 => "0100000001001011",
5787 => "0100000001001011",5788 => "0100001011101111",
5789 => "0100001011110000",5790 => "0100001011110001",
5791 => "0100001011110010",5792 => "0100001011110011",
5793 => "0100001011110100",5794 => "0100001011110101",
5795 => "0100001011110101",5796 => "0100001011110110",
5797 => "0100001011110111",5798 => "0100000001001100",
5799 => "0100001011111001",5800 => "0100001011111010",
5801 => "0100001011111011",5802 => "0100001011111100",
5803 => "0100001011111100",5804 => "0100001011111101",
5805 => "0100001011111110",5806 => "0100001011111111",
5807 => "0100001100000000",5808 => "0100001100000001",
5809 => "0100000001001101",5810 => "0100001100000011",
5811 => "0100001100000011",5812 => "0100001100000100",
5813 => "0100001100000101",5814 => "0100001100000110",
5815 => "0100001100000111",5816 => "0100001100001000",
5817 => "0100001100001001",5818 => "0100001100001010",
5819 => "0100001100001010",5820 => "0100001100001011",
5821 => "0100000001001110",5822 => "0100001100001101",
5823 => "0100001100001110",5824 => "0100001100001111",
5825 => "0100001100010000",5826 => "0100001100010001",
5827 => "0100001100010001",5828 => "0100001100010010",
5829 => "0100001100010011",5830 => "0100001100010100",
5831 => "0100001100010101",5832 => "0100000001001111",
5833 => "0100001100010111",5834 => "0100001100011000",
5835 => "0100001100011001",5836 => "0100001100011001",
5837 => "0100001100011010",5838 => "0100001100011011",
5839 => "0100001100011100",5840 => "0100001100011101",
5841 => "0100001100011110",5842 => "0100001100011111",
5843 => "0100000000001000",5844 => "0100000000001000",
5845 => "0100001100100001",5846 => "0100001100100010",
5847 => "0100001100100011",5848 => "0100001100100100",
5849 => "0100001100100101",5850 => "0100001100100110",
5851 => "0100001100100111",5852 => "0100001100100111",
5853 => "0100001100101000",5854 => "0100001100101001",
5855 => "0100000001010001",5856 => "0100001100101011",
5857 => "0100001100101100",5858 => "0100001100101101",
5859 => "0100001100101110",5860 => "0100001100101111",
5861 => "0100001100101111",5862 => "0100001100110000",
5863 => "0100001100110001",5864 => "0100001100110010",
5865 => "0100001100110011",5866 => "0100000001010010",
5867 => "0100001100110101",5868 => "0100001100110110",
5869 => "0100001100110110",5870 => "0100001100110111",
5871 => "0100001100111000",5872 => "0100001100111001",
5873 => "0100001100111010",5874 => "0100001100111011",
5875 => "0100001100111100",5876 => "0100001100111101",
5877 => "0100000001010011",5878 => "0100000001010011",
5879 => "0100001100111111",5880 => "0100001101000000",
5881 => "0100001101000001",5882 => "0100001101000010",
5883 => "0100001101000011",5884 => "0100001101000100",
5885 => "0100001101000101",5886 => "0100001101000101",
5887 => "0100001101000110",5888 => "0100001101000111",
5889 => "0100000001010100",5890 => "0100001101001001",
5891 => "0100001101001010",5892 => "0100001101001011",
5893 => "0100001101001100",5894 => "0100001101001101",
5895 => "0100001101001101",5896 => "0100001101001110",
5897 => "0100001101001111",5898 => "0100001101010000",
5899 => "0100001101010001",5900 => "0100000001010101",
5901 => "0100001101010011",5902 => "0100001101010100",
5903 => "0100001101010101",5904 => "0100001101010101",
5905 => "0100001101010110",5906 => "0100001101010111",
5907 => "0100001101011000",5908 => "0100001101011001",
5909 => "0100001101011010",5910 => "0100001101011011",
5911 => "0100000001010110",5912 => "0100000001010110",
5913 => "0100001101011101",5914 => "0100001101011110",
5915 => "0100001101011111",5916 => "0100001101100000",
5917 => "0100001101100001",5918 => "0100001101100010",
5919 => "0100001101100011",5920 => "0100001101100100",
5921 => "0100001101100100",5922 => "0100001101100101",
5923 => "0100000001010111",5924 => "0100001101100111",
5925 => "0100001101101000",5926 => "0100001101101001",
5927 => "0100001101101010",5928 => "0100001101101011",
5929 => "0100001101101100",5930 => "0100001101101100",
5931 => "0100001101101101",5932 => "0100001101101110",
5933 => "0100001101101111",5934 => "0100000001011000",
5935 => "0100001101110001",5936 => "0100001101110010",
5937 => "0100001101110011",5938 => "0100001101110100",
5939 => "0100001101110100",5940 => "0100001101110101",
5941 => "0100001101110110",5942 => "0100001101110111",
5943 => "0100001101111000",5944 => "0100001101111001",
5945 => "0100000001011001",5946 => "0100001101111011",
5947 => "0100001101111100",5948 => "0100001101111100",
5949 => "0100001101111101",5950 => "0100001101111110",
5951 => "0100001101111111",5952 => "0100001110000000",
5953 => "0100001110000001",5954 => "0100001110000010",
5955 => "0100001110000011",5956 => "0100000000001001",
5957 => "0100000000001001",5958 => "0100001110000101",
5959 => "0100001110000110",5960 => "0100001110000111",
5961 => "0100001110001000",5962 => "0100001110001001",
5963 => "0100001110001010",5964 => "0100001110001011",
5965 => "0100001110001100",5966 => "0100001110001100",
5967 => "0100001110001101",5968 => "0100000001011011",
5969 => "0100001110001111",5970 => "0100001110010000",
5971 => "0100001110010001",5972 => "0100001110010010",
5973 => "0100001110010011",5974 => "0100001110010100",
5975 => "0100001110010100",5976 => "0100001110010101",
5977 => "0100001110010110",5978 => "0100001110010111",
5979 => "0100000001011100",5980 => "0100001110011001",
5981 => "0100001110011010",5982 => "0100001110011011",
5983 => "0100001110011100",5984 => "0100001110011100",
5985 => "0100001110011101",5986 => "0100001110011110",
5987 => "0100001110011111",5988 => "0100001110100000",
5989 => "0100001110100001",5990 => "0100000001011101",
5991 => "0100001110100011",5992 => "0100001110100100",
5993 => "0100001110100101",5994 => "0100001110100101",
5995 => "0100001110100110",5996 => "0100001110100111",
5997 => "0100001110101000",5998 => "0100001110101001",
5999 => "0100001110101010",6000 => "0100001110101011",
6001 => "0100000001011110",6002 => "0100001110101101",
6003 => "0100001110101101",6004 => "0100001110101110",
6005 => "0100001110101111",6006 => "0100001110110000",
6007 => "0100001110110001",6008 => "0100001110110010",
6009 => "0100001110110011",6010 => "0100001110110100",
6011 => "0100001110110101",6012 => "0100000001011111",
6013 => "0100000001011111",6014 => "0100001110110111",
6015 => "0100001110111000",6016 => "0100001110111001",
6017 => "0100001110111010",6018 => "0100001110111011",
6019 => "0100001110111100",6020 => "0100001110111101",
6021 => "0100001110111110",6022 => "0100001110111110",
6023 => "0100001110111111",6024 => "0100000001100000",
6025 => "0100001111000001",6026 => "0100001111000010",
6027 => "0100001111000011",6028 => "0100001111000100",
6029 => "0100001111000101",6030 => "0100001111000110",
6031 => "0100001111000111",6032 => "0100001111000111",
6033 => "0100001111001000",6034 => "0100001111001001",
6035 => "0100000001100001",6036 => "0100001111001011",
6037 => "0100001111001100",6038 => "0100001111001101",
6039 => "0100001111001110",6040 => "0100001111001111",
6041 => "0100001111010000",6042 => "0100001111010000",
6043 => "0100001111010001",6044 => "0100001111010010",
6045 => "0100001111010011",6046 => "0100000001100010",
6047 => "0100001111010101",6048 => "0100001111010110",
6049 => "0100001111010111",6050 => "0100001111011000",
6051 => "0100001111011000",6052 => "0100001111011001",
6053 => "0100001111011010",6054 => "0100001111011011",
6055 => "0100001111011100",6056 => "0100001111011101",
6057 => "0100000001100011",6058 => "0100001111011111",
6059 => "0100001111100000",6060 => "0100001111100001",
6061 => "0100001111100001",6062 => "0100001111100010",
6063 => "0100001111100011",6064 => "0100001111100100",
6065 => "0100001111100101",6066 => "0100001111100110",
6067 => "0100001111100111",6068 => "0100100000000000",
6069 => "0100100000000001",6070 => "0100100000000010",
6071 => "0100100000000010",6072 => "0100100000000011",
6073 => "0100100000000100",6074 => "0100100000000101",
6075 => "0100100000000110",6076 => "0100100000000111",
6077 => "0100100000001000",6078 => "0100100000001001",
6079 => "0100100000000001",6080 => "0100100000001011",
6081 => "0100100000001011",6082 => "0100100000001100",
6083 => "0100100000001101",6084 => "0100100000001110",
6085 => "0100100000001111",6086 => "0100100000010000",
6087 => "0100100000010001",6088 => "0100100000010010",
6089 => "0100100000010011",6090 => "0100100000000010",
6091 => "0100100000010101",6092 => "0100100000010101",
6093 => "0100100000010110",6094 => "0100100000010111",
6095 => "0100100000011000",6096 => "0100100000011001",
6097 => "0100100000011010",6098 => "0100100000011011",
6099 => "0100100000011100",6100 => "0100100000011101",
6101 => "0100100000000011",6102 => "0100100000000011",
6103 => "0100100000011111",6104 => "0100100000100000",
6105 => "0100100000100001",6106 => "0100100000100010",
6107 => "0100100000100011",6108 => "0100100000100100",
6109 => "0100100000100101",6110 => "0100100000100110",
6111 => "0100100000100111",6112 => "0100100000100111",
6113 => "0100100000000100",6114 => "0100100000101001",
6115 => "0100100000101010",6116 => "0100100000101011",
6117 => "0100100000101100",6118 => "0100100000101101",
6119 => "0100100000101110",6120 => "0100100000101111",
6121 => "0100100000110000",6122 => "0100100000110001",
6123 => "0100100000110001",6124 => "0100100000000101",
6125 => "0100100000110011",6126 => "0100100000110100",
6127 => "0100100000110101",6128 => "0100100000110110",
6129 => "0100100000110111",6130 => "0100100000111000",
6131 => "0100100000111001",6132 => "0100100000111010",
6133 => "0100100000111010",6134 => "0100100000111011",
6135 => "0100100000000110",6136 => "0100100000111101",
6137 => "0100100000111110",6138 => "0100100000111111",
6139 => "0100100001000000",6140 => "0100100001000001",
6141 => "0100100001000010",6142 => "0100100001000011",
6143 => "0100100001000100",6144 => "0000000000000000",
6145 => "0000000000000000",6146 => "0000000000000000",
6147 => "0000000000000000",6148 => "0000000000000000",
6149 => "0000000000000000",6150 => "0000000000000000",
6151 => "0000000000000000",6152 => "0000000000000000",
6153 => "0000000000000000",6154 => "0000000000000000",
6155 => "0000000000000000",6156 => "0000000000000000",
6157 => "0000000000000000",6158 => "0000000000000000",
6159 => "0000000000000000",6160 => "0000000000000000",
6161 => "0000000000000000",6162 => "0000000000000000",
6163 => "0000000000000000",6164 => "0000000000000000",
6165 => "0000000000000000",6166 => "0000000000000000",
6167 => "0000000000000000",6168 => "0000000000000000",
6169 => "0000000000000000",6170 => "0000000000000000",
6171 => "0000000000000000",6172 => "0000000000000000",
6173 => "0000000000000000",6174 => "0000000000000000",
6175 => "0000000000000000",6176 => "0000000000000000",
6177 => "0000000000000000",6178 => "0000000000000000",
6179 => "0000000000000000",6180 => "0000000000000000",
6181 => "0000000000000000",6182 => "0000000000000000",
6183 => "0000000000000000",6184 => "0000000000000000",
6185 => "0000000000000000",6186 => "0000000000000000",
6187 => "0000000000000000",6188 => "0000000000000000",
6189 => "0000000000000000",6190 => "0000000000000000",
6191 => "0000000000000000",6192 => "0000000000000000",
6193 => "0000000000000000",6194 => "0000000000000000",
6195 => "0000000000000000",6196 => "0000000000000000",
6197 => "0000000000000000",6198 => "0000000000000000",
6199 => "0000000000000000",6200 => "0000000000000000",
6201 => "0000000000000000",6202 => "0000000000000000",
6203 => "0000000000000000",6204 => "0000000000000000",
6205 => "0000000000000000",6206 => "0000000000000000",
6207 => "0000000000000000",6208 => "0000000000000000",
6209 => "0000000000000000",6210 => "0000000000000000",
6211 => "0000000000000000",6212 => "0000000000000000",
6213 => "0000000000000000",6214 => "0000000000000000",
6215 => "0000000000000000",6216 => "0000000000000000",
6217 => "0000000000000000",6218 => "0000000000000000",
6219 => "0000000000000000",6220 => "0000000000000000",
6221 => "0000000000000000",6222 => "0000000000000000",
6223 => "0000000000000000",6224 => "0000000000000000",
6225 => "0000000000000000",6226 => "0000000000000000",
6227 => "0000000000000000",6228 => "0000000000000000",
6229 => "0000000000000000",6230 => "0000000000000000",
6231 => "0000000000000000",6232 => "0000000000000000",
6233 => "0000000000000000",6234 => "0000000000000000",
6235 => "0000000000000000",6236 => "0000000000000000",
6237 => "0000000000000000",6238 => "0000000000000000",
6239 => "0000000000000000",6240 => "0000000000000000",
6241 => "0000000000000000",6242 => "0000000000000000",
6243 => "0000000000000000",6244 => "0000000000000000",
6245 => "0000000000000000",6246 => "0000000000000000",
6247 => "0000000000000000",6248 => "0000000000000000",
6249 => "0000000000000000",6250 => "0000000000000000",
6251 => "0000000000000000",6252 => "0000000000000000",
6253 => "0000000000000000",6254 => "0000000000000000",
6255 => "0000000000000000",6256 => "0000000000000000",
6257 => "0000000000000000",6258 => "0000000000000000",
6259 => "0000000000000000",6260 => "0000000000000000",
6261 => "0000000000000000",6262 => "0000000000000000",
6263 => "0000000000000000",6264 => "0000000000000000",
6265 => "0000000000000000",6266 => "0000000000000000",
6267 => "0000000000000000",6268 => "0000000000000000",
6269 => "0000000000000000",6270 => "0000000000000000",
6271 => "0000000000000000",6272 => "0000000000000000",
6273 => "0000000000000000",6274 => "0000000000000000",
6275 => "0000000000000000",6276 => "0000000000000000",
6277 => "0000000000000000",6278 => "0000000000000000",
6279 => "0000000000000000",6280 => "0000000000000000",
6281 => "0000000000000000",6282 => "0000000000000000",
6283 => "0000000000000000",6284 => "0000000000000000",
6285 => "0000000000000000",6286 => "0000000000000000",
6287 => "0000000000000000",6288 => "0000000000000000",
6289 => "0000000000000000",6290 => "0000000000000000",
6291 => "0000000000000000",6292 => "0000000000000000",
6293 => "0000000000000000",6294 => "0000000000000000",
6295 => "0000000000000000",6296 => "0000000000000000",
6297 => "0000000000000000",6298 => "0000000000000000",
6299 => "0000000000000000",6300 => "0000000000000000",
6301 => "0000000000000000",6302 => "0000000000000000",
6303 => "0000000000000000",6304 => "0000000000000000",
6305 => "0000000000000000",6306 => "0000000000000000",
6307 => "0000000000000000",6308 => "0000000000000000",
6309 => "0000000000000000",6310 => "0000000000000000",
6311 => "0000000000000000",6312 => "0000000000000000",
6313 => "0000000000000000",6314 => "0000000000000000",
6315 => "0000000000000000",6316 => "0000000000000000",
6317 => "0000000000000000",6318 => "0000000000000000",
6319 => "0000000000000000",6320 => "0000000000000000",
6321 => "0000000000000000",6322 => "0000000000000000",
6323 => "0000000000000000",6324 => "0000000000000000",
6325 => "0000000000000000",6326 => "0000000000000000",
6327 => "0000000000000000",6328 => "0000000000000000",
6329 => "0000000000000000",6330 => "0000000000000000",
6331 => "0000000000000000",6332 => "0000000000000000",
6333 => "0000000000000000",6334 => "0000000000000000",
6335 => "0000000000000000",6336 => "0000000000000000",
6337 => "0000000000000000",6338 => "0000000000000000",
6339 => "0000000000000000",6340 => "0000000000000000",
6341 => "0000000000000000",6342 => "0000000000000000",
6343 => "0000000000000000",6344 => "0000000000000000",
6345 => "0000000000000000",6346 => "0000000000000000",
6347 => "0000000000000000",6348 => "0000000000000000",
6349 => "0000000000000000",6350 => "0000000000000000",
6351 => "0000000000000000",6352 => "0000000000000000",
6353 => "0000000000000000",6354 => "0000000000000000",
6355 => "0000000000000000",6356 => "0000000000000000",
6357 => "0000000000000000",6358 => "0000000000000000",
6359 => "0000000000000000",6360 => "0000000000000000",
6361 => "0000000000000000",6362 => "0000000000000000",
6363 => "0000000000000000",6364 => "0000000000000000",
6365 => "0000000000000000",6366 => "0000000000000000",
6367 => "0000000000000000",6368 => "0000000000000000",
6369 => "0000000000000000",6370 => "0000000000000000",
6371 => "0000000000000000",6372 => "0000000000000000",
6373 => "0000000000000000",6374 => "0000000000000000",
6375 => "0000000000000000",6376 => "0000000000000000",
6377 => "0000000000000000",6378 => "0000000000000000",
6379 => "0000000000000000",6380 => "0000000000000000",
6381 => "0000000000000000",6382 => "0000000000000000",
6383 => "0000000000000000",6384 => "0000000000000000",
6385 => "0000000000000000",6386 => "0000000000000000",
6387 => "0000000000000000",6388 => "0000000000000000",
6389 => "0000000000000000",6390 => "0000000000000000",
6391 => "0000000000000000",6392 => "0000000000000000",
6393 => "0000000000000000",6394 => "0000000000000000",
6395 => "0000000000000000",6396 => "0000000000000000",
6397 => "0000000000000000",6398 => "0000000000000000",
6399 => "0000000000000000",6400 => "0000000000000000",
6401 => "0000000000000000",6402 => "0000000000000000",
6403 => "0000000000000000",6404 => "0000000000000000",
6405 => "0000000000000000",6406 => "0000000000000000",
6407 => "0000000000000000",6408 => "0000000000000000",
6409 => "0000000000000000",6410 => "0000000000000000",
6411 => "0000000000000000",6412 => "0000000000000000",
6413 => "0000000000000000",6414 => "0000000000000000",
6415 => "0000000000000000",6416 => "0000000000000000",
6417 => "0000000000000000",6418 => "0000000000000000",
6419 => "0000000000000000",6420 => "0000000000000000",
6421 => "0000000000000000",6422 => "0000000000000000",
6423 => "0000000000000000",6424 => "0000000000000000",
6425 => "0000000000000000",6426 => "0000000000000000",
6427 => "0000000000000000",6428 => "0000000000000000",
6429 => "0000000000000000",6430 => "0000000000000000",
6431 => "0000000000000000",6432 => "0000000000000000",
6433 => "0000000000000000",6434 => "0000000000000000",
6435 => "0000000000000000",6436 => "0000000000000000",
6437 => "0000000000000000",6438 => "0000000000000000",
6439 => "0000000000000000",6440 => "0000000000000000",
6441 => "0000000000000000",6442 => "0000000000000000",
6443 => "0000000000000000",6444 => "0000000000000000",
6445 => "0000000000000000",6446 => "0000000000000000",
6447 => "0000000000000000",6448 => "0000000000000000",
6449 => "0000000000000000",6450 => "0000000000000000",
6451 => "0000000000000000",6452 => "0000000000000000",
6453 => "0000000000000000",6454 => "0000000000000000",
6455 => "0000000000000000",6456 => "0000000000000000",
6457 => "0000000000000000",6458 => "0000000000000000",
6459 => "0000000000000000",6460 => "0000000000000000",
6461 => "0000000000000000",6462 => "0000000000000000",
6463 => "0000000000000000",6464 => "0000000000000000",
6465 => "0000000000000000",6466 => "0000000000000000",
6467 => "0000000000000000",6468 => "0000000000000000",
6469 => "0000000000000000",6470 => "0000000000000000",
6471 => "0000000000000000",6472 => "0000000000000000",
6473 => "0000000000000000",6474 => "0000000000000000",
6475 => "0000000000000000",6476 => "0000000000000000",
6477 => "0000000000000000",6478 => "0000000000000000",
6479 => "0000000000000000",6480 => "0000000000000000",
6481 => "0000000000000000",6482 => "0000000000000000",
6483 => "0000000000000000",6484 => "0000000000000000",
6485 => "0000000000000000",6486 => "0000000000000000",
6487 => "0000000000000000",6488 => "0000000000000000",
6489 => "0000000000000000",6490 => "0000000000000000",
6491 => "0000000000000000",6492 => "0000000000000000",
6493 => "0000000000000000",6494 => "0000000000000000",
6495 => "0000000000000000",6496 => "0000000000000000",
6497 => "0000000000000000",6498 => "0000000000000000",
6499 => "0000000000000000",6500 => "0000000000000000",
6501 => "0000000000000000",6502 => "0000000000000000",
6503 => "0000000000000000",6504 => "0000000000000000",
6505 => "0000000000000000",6506 => "0000000000000000",
6507 => "0000000000000000",6508 => "0000000000000000",
6509 => "0000000000000000",6510 => "0000000000000000",
6511 => "0000000000000000",6512 => "0000000000000000",
6513 => "0000000000000000",6514 => "0000000000000000",
6515 => "0000000000000000",6516 => "0000000000000000",
6517 => "0000000000000000",6518 => "0000000000000000",
6519 => "0000000000000000",6520 => "0000000000000000",
6521 => "0000000000000000",6522 => "0000000000000000",
6523 => "0000000000000000",6524 => "0000000000000000",
6525 => "0000000000000000",6526 => "0000000000000000",
6527 => "0000000000000000",6528 => "0000000000000000",
6529 => "0000000000000000",6530 => "0000000000000000",
6531 => "0000000000000000",6532 => "0000000000000000",
6533 => "0000000000000000",6534 => "0000000000000000",
6535 => "0000000000000000",6536 => "0000000000000000",
6537 => "0000000000000000",6538 => "0000000000000000",
6539 => "0000000000000000",6540 => "0000000000000000",
6541 => "0000000000000000",6542 => "0000000000000000",
6543 => "0000000000000000",6544 => "0000000000000000",
6545 => "0000000000000000",6546 => "0000000000000000",
6547 => "0000000000000000",6548 => "0000000000000000",
6549 => "0000000000000000",6550 => "0000000000000000",
6551 => "0000000000000000",6552 => "0000000000000000",
6553 => "0000000000000000",6554 => "0000000000000000",
6555 => "0000000000000000",6556 => "0000000000000000",
6557 => "0000000000000000",6558 => "0000000000000000",
6559 => "0000000000000000",6560 => "0000000000000000",
6561 => "0000000000000000",6562 => "0000000000000000",
6563 => "0000000000000000",6564 => "0000000000000000",
6565 => "0000000000000000",6566 => "0000000000000000",
6567 => "0000000000000000",6568 => "0000000000000000",
6569 => "0000000000000000",6570 => "0000000000000000",
6571 => "0000000000000000",6572 => "0000000000000000",
6573 => "0000000000000000",6574 => "0000000000000000",
6575 => "0000000000000000",6576 => "0000000000000000",
6577 => "0000000000000000",6578 => "0000000000000000",
6579 => "0000000000000000",6580 => "0000000000000000",
6581 => "0000000000000000",6582 => "0000000000000000",
6583 => "0000000000000000",6584 => "0000000000000000",
6585 => "0000000000000000",6586 => "0000000000000000",
6587 => "0000000000000000",6588 => "0000000000000000",
6589 => "0000000000000000",6590 => "0000000000000000",
6591 => "0000000000000000",6592 => "0000000000000000",
6593 => "0000000000000000",6594 => "0000000000000000",
6595 => "0000000000000000",6596 => "0000000000000000",
6597 => "0000000000000000",6598 => "0000000000000000",
6599 => "0000000000000000",6600 => "0000000000000000",
6601 => "0000000000000000",6602 => "0000000000000000",
6603 => "0000000000000000",6604 => "0000000000000000",
6605 => "0000000000000000",6606 => "0000000000000000",
6607 => "0000000000000000",6608 => "0000000000000000",
6609 => "0000000000000000",6610 => "0000000000000000",
6611 => "0000000000000000",6612 => "0000000000000000",
6613 => "0000000000000000",6614 => "0000000000000000",
6615 => "0000000000000000",6616 => "0000000000000000",
6617 => "0000000000000000",6618 => "0000000000000000",
6619 => "0000000000000000",6620 => "0000000000000000",
6621 => "0000000000000000",6622 => "0000000000000000",
6623 => "0000000000000000",6624 => "0000000000000000",
6625 => "0000000000000000",6626 => "0000000000000000",
6627 => "0000000000000000",6628 => "0000000000000000",
6629 => "0000000000000000",6630 => "0000000000000000",
6631 => "0000000000000000",6632 => "0000000000000000",
6633 => "0000000000000000",6634 => "0000000000000000",
6635 => "0000000000000000",6636 => "0000000000000000",
6637 => "0000000000000000",6638 => "0000000000000000",
6639 => "0000000000000000",6640 => "0000000000000000",
6641 => "0000000000000000",6642 => "0000000000000000",
6643 => "0000000000000000",6644 => "0000000000000000",
6645 => "0000000000000000",6646 => "0000000000000000",
6647 => "0000000000000000",6648 => "0000000000000000",
6649 => "0000000000000000",6650 => "0000000000000000",
6651 => "0000000000000000",6652 => "0000000000000000",
6653 => "0000000000000000",6654 => "0000000000000000",
6655 => "0000000000000000",6656 => "0000000000000000",
6657 => "0000000000000000",6658 => "0000000000000000",
6659 => "0000000000000000",6660 => "0000000000000000",
6661 => "0000000000000000",6662 => "0000000000000000",
6663 => "0000000000000000",6664 => "0000000000000000",
6665 => "0000000000000000",6666 => "0000000000000000",
6667 => "0000000000000000",6668 => "0000000000000000",
6669 => "0000000000000000",6670 => "0000000000000000",
6671 => "0000000000000000",6672 => "0000000000000000",
6673 => "0000000000000000",6674 => "0000000000000000",
6675 => "0000000000000000",6676 => "0000000000000000",
6677 => "0000000000000000",6678 => "0000000000000000",
6679 => "0000000000000000",6680 => "0000000000000000",
6681 => "0000000000000000",6682 => "0000000000000000",
6683 => "0000000000000000",6684 => "0000000000000000",
6685 => "0000000000000000",6686 => "0000000000000000",
6687 => "0000000000000000",6688 => "0000000000000000",
6689 => "0000000000000000",6690 => "0000000000000000",
6691 => "0000000000000000",6692 => "0000000000000000",
6693 => "0000000000000000",6694 => "0000000000000000",
6695 => "0000000000000000",6696 => "0000000000000000",
6697 => "0000000000000000",6698 => "0000000000000000",
6699 => "0000000000000000",6700 => "0000000000000000",
6701 => "0000000000000000",6702 => "0000000000000000",
6703 => "0000000000000000",6704 => "0000000000000000",
6705 => "0000000000000000",6706 => "0000000000000000",
6707 => "0000000000000000",6708 => "0000000000000000",
6709 => "0000000000000000",6710 => "0000000000000000",
6711 => "0000000000000000",6712 => "0000000000000000",
6713 => "0000000000000000",6714 => "0000000000000000",
6715 => "0000000000000000",6716 => "0000000000000000",
6717 => "0000000000000000",6718 => "0000000000000000",
6719 => "0000000000000000",6720 => "0000000000000000",
6721 => "0000000000000000",6722 => "0000000000000000",
6723 => "0000000000000000",6724 => "0000000000000000",
6725 => "0000000000000000",6726 => "0000000000000000",
6727 => "0000000000000000",6728 => "0000000000000000",
6729 => "0000000000000000",6730 => "0000000000000000",
6731 => "0000000000000000",6732 => "0000000000000000",
6733 => "0000000000000000",6734 => "0000000000000000",
6735 => "0000000000000000",6736 => "0000000000000000",
6737 => "0000000000000000",6738 => "0000000000000000",
6739 => "0000000000000000",6740 => "0000000000000000",
6741 => "0000000000000000",6742 => "0000000000000000",
6743 => "0000000000000000",6744 => "0000000000000000",
6745 => "0000000000000000",6746 => "0000000000000000",
6747 => "0000000000000000",6748 => "0000000000000000",
6749 => "0000000000000000",6750 => "0000000000000000",
6751 => "0000000000000000",6752 => "0000000000000000",
6753 => "0000000000000000",6754 => "0000000000000000",
6755 => "0000000000000000",6756 => "0000000000000000",
6757 => "0000000000000000",6758 => "0000000000000000",
6759 => "0000000000000000",6760 => "0000000000000000",
6761 => "0000000000000000",6762 => "0000000000000000",
6763 => "0000000000000000",6764 => "0000000000000000",
6765 => "0000000000000000",6766 => "0000000000000000",
6767 => "0000000000000000",6768 => "0000000000000000",
6769 => "0000000000000000",6770 => "0000000000000000",
6771 => "0000000000000000",6772 => "0000000000000000",
6773 => "0000000000000000",6774 => "0000000000000000",
6775 => "0000000000000000",6776 => "0000000000000000",
6777 => "0000000000000000",6778 => "0000000000000000",
6779 => "0000000000000000",6780 => "0000000000000000",
6781 => "0000000000000000",6782 => "0000000000000000",
6783 => "0000000000000000",6784 => "0000000000000000",
6785 => "0000000000000000",6786 => "0000000000000000",
6787 => "0000000000000000",6788 => "0000000000000000",
6789 => "0000000000000000",6790 => "0000000000000000",
6791 => "0000000000000000",6792 => "0000000000000000",
6793 => "0000000000000000",6794 => "0000000000000000",
6795 => "0000000000000000",6796 => "0000000000000000",
6797 => "0000000000000000",6798 => "0000000000000000",
6799 => "0000000000000000",6800 => "0000000000000000",
6801 => "0000000000000000",6802 => "0000000000000000",
6803 => "0000000000000000",6804 => "0000000000000000",
6805 => "0000000000000000",6806 => "0000000000000000",
6807 => "0000000000000000",6808 => "0000000000000000",
6809 => "0000000000000000",6810 => "0000000000000000",
6811 => "0000000000000000",6812 => "0000000000000000",
6813 => "0000000000000000",6814 => "0000000000000000",
6815 => "0000000000000000",6816 => "0000000000000000",
6817 => "0000000000000000",6818 => "0000000000000000",
6819 => "0000000000000000",6820 => "0000000000000000",
6821 => "0000000000000000",6822 => "0000000000000000",
6823 => "0000000000000000",6824 => "0000000000000000",
6825 => "0000000000000000",6826 => "0000000000000000",
6827 => "0000000000000000",6828 => "0000000000000000",
6829 => "0000000000000000",6830 => "0000000000000000",
6831 => "0000000000000000",6832 => "0000000000000000",
6833 => "0000000000000000",6834 => "0000000000000000",
6835 => "0000000000000000",6836 => "0000000000000000",
6837 => "0000000000000000",6838 => "0000000000000000",
6839 => "0000000000000000",6840 => "0000000000000000",
6841 => "0000000000000000",6842 => "0000000000000000",
6843 => "0000000000000000",6844 => "0000000000000000",
6845 => "0000000000000000",6846 => "0000000000000000",
6847 => "0000000000000000",6848 => "0000000000000000",
6849 => "0000000000000000",6850 => "0000000000000000",
6851 => "0000000000000000",6852 => "0000000000000000",
6853 => "0000000000000000",6854 => "0000000000000000",
6855 => "0000000000000000",6856 => "0000000000000000",
6857 => "0000000000000000",6858 => "0000000000000000",
6859 => "0000000000000000",6860 => "0000000000000000",
6861 => "0000000000000000",6862 => "0000000000000000",
6863 => "0000000000000000",6864 => "0000000000000000",
6865 => "0000000000000000",6866 => "0000000000000000",
6867 => "0000000000000000",6868 => "0000000000000000",
6869 => "0000000000000000",6870 => "0000000000000000",
6871 => "0000000000000000",6872 => "0000000000000000",
6873 => "0000000000000000",6874 => "0000000000000000",
6875 => "0000000000000000",6876 => "0000000000000000",
6877 => "0000000000000000",6878 => "0000000000000000",
6879 => "0000000000000000",6880 => "0000000000000000",
6881 => "0000000000000000",6882 => "0000000000000000",
6883 => "0000000000000000",6884 => "0000000000000000",
6885 => "0000000000000000",6886 => "0000000000000000",
6887 => "0000000000000000",6888 => "0000000000000000",
6889 => "0000000000000000",6890 => "0000000000000000",
6891 => "0000000000000000",6892 => "0000000000000000",
6893 => "0000000000000000",6894 => "0000000000000000",
6895 => "0000000000000000",6896 => "0000000000000000",
6897 => "0000000000000000",6898 => "0000000000000000",
6899 => "0000000000000000",6900 => "0000000000000000",
6901 => "0000000000000000",6902 => "0000000000000000",
6903 => "0000000000000000",6904 => "0000000000000000",
6905 => "0000000000000000",6906 => "0000000000000000",
6907 => "0000000000000000",6908 => "0000000000000000",
6909 => "0000000000000000",6910 => "0000000000000000",
6911 => "0000000000000000",6912 => "0000000000000000",
6913 => "0000000000000000",6914 => "0000000000000000",
6915 => "0000000000000000",6916 => "0000000000000000",
6917 => "0000000000000000",6918 => "0000000000000000",
6919 => "0000000000000000",6920 => "0000000000000000",
6921 => "0000000000000000",6922 => "0000000000000000",
6923 => "0000000000000000",6924 => "0000000000000000",
6925 => "0000000000000000",6926 => "0000000000000000",
6927 => "0000000000000000",6928 => "0000000000000000",
6929 => "0000000000000000",6930 => "0000000000000000",
6931 => "0000000000000000",6932 => "0000000000000000",
6933 => "0000000000000000",6934 => "0000000000000000",
6935 => "0000000000000000",6936 => "0000000000000000",
6937 => "0000000000000000",6938 => "0000000000000000",
6939 => "0000000000000000",6940 => "0000000000000000",
6941 => "0000000000000000",6942 => "0000000000000000",
6943 => "0000000000000000",6944 => "0000000000000000",
6945 => "0000000000000000",6946 => "0000000000000000",
6947 => "0000000000000000",6948 => "0000000000000000",
6949 => "0000000000000000",6950 => "0000000000000000",
6951 => "0000000000000000",6952 => "0000000000000000",
6953 => "0000000000000000",6954 => "0000000000000000",
6955 => "0000000000000000",6956 => "0000000000000000",
6957 => "0000000000000000",6958 => "0000000000000000",
6959 => "0000000000000000",6960 => "0000000000000000",
6961 => "0000000000000000",6962 => "0000000000000000",
6963 => "0000000000000000",6964 => "0000000000000000",
6965 => "0000000000000000",6966 => "0000000000000000",
6967 => "0000000000000000",6968 => "0000000000000000",
6969 => "0000000000000000",6970 => "0000000000000000",
6971 => "0000000000000000",6972 => "0000000000000000",
6973 => "0000000000000000",6974 => "0000000000000000",
6975 => "0000000000000000",6976 => "0000000000000000",
6977 => "0000000000000000",6978 => "0000000000000000",
6979 => "0000000000000000",6980 => "0000000000000000",
6981 => "0000000000000000",6982 => "0000000000000000",
6983 => "0000000000000000",6984 => "0000000000000000",
6985 => "0000000000000000",6986 => "0000000000000000",
6987 => "0000000000000000",6988 => "0000000000000000",
6989 => "0000000000000000",6990 => "0000000000000000",
6991 => "0000000000000000",6992 => "0000000000000000",
6993 => "0000000000000000",6994 => "0000000000000000",
6995 => "0000000000000000",6996 => "0000000000000000",
6997 => "0000000000000000",6998 => "0000000000000000",
6999 => "0000000000000000",7000 => "0000000000000000",
7001 => "0000000000000000",7002 => "0000000000000000",
7003 => "0000000000000000",7004 => "0000000000000000",
7005 => "0000000000000000",7006 => "0000000000000000",
7007 => "0000000000000000",7008 => "0000000000000000",
7009 => "0000000000000000",7010 => "0000000000000000",
7011 => "0000000000000000",7012 => "0000000000000000",
7013 => "0000000000000000",7014 => "0000000000000000",
7015 => "0000000000000000",7016 => "0000000000000000",
7017 => "0000000000000000",7018 => "0000000000000000",
7019 => "0000000000000000",7020 => "0000000000000000",
7021 => "0000000000000000",7022 => "0000000000000000",
7023 => "0000000000000000",7024 => "0000000000000000",
7025 => "0000000000000000",7026 => "0000000000000000",
7027 => "0000000000000000",7028 => "0000000000000000",
7029 => "0000000000000000",7030 => "0000000000000000",
7031 => "0000000000000000",7032 => "0000000000000000",
7033 => "0000000000000000",7034 => "0000000000000000",
7035 => "0000000000000000",7036 => "0000000000000000",
7037 => "0000000000000000",7038 => "0000000000000000",
7039 => "0000000000000000",7040 => "0000000000000000",
7041 => "0000000000000000",7042 => "0000000000000000",
7043 => "0000000000000000",7044 => "0000000000000000",
7045 => "0000000000000000",7046 => "0000000000000000",
7047 => "0000000000000000",7048 => "0000000000000000",
7049 => "0000000000000000",7050 => "0000000000000000",
7051 => "0000000000000000",7052 => "0000000000000000",
7053 => "0000000000000000",7054 => "0000000000000000",
7055 => "0000000000000000",7056 => "0000000000000000",
7057 => "0000000000000000",7058 => "0000000000000000",
7059 => "0000000000000000",7060 => "0000000000000000",
7061 => "0000000000000000",7062 => "0000000000000000",
7063 => "0000000000000000",7064 => "0000000000000000",
7065 => "0000000000000000",7066 => "0000000000000000",
7067 => "0000000000000000",7068 => "0000000000000000",
7069 => "0000000000000000",7070 => "0000000000000000",
7071 => "0000000000000000",7072 => "0000000000000000",
7073 => "0000000000000000",7074 => "0000000000000000",
7075 => "0000000000000000",7076 => "0000000000000000",
7077 => "0000000000000000",7078 => "0000000000000000",
7079 => "0000000000000000",7080 => "0000000000000000",
7081 => "0000000000000000",7082 => "0000000000000000",
7083 => "0000000000000000",7084 => "0000000000000000",
7085 => "0000000000000000",7086 => "0000000000000000",
7087 => "0000000000000000",7088 => "0000000000000000",
7089 => "0000000000000000",7090 => "0000000000000000",
7091 => "0000000000000000",7092 => "0000000000000000",
7093 => "0000000000000000",7094 => "0000000000000000",
7095 => "0000000000000000",7096 => "0000000000000000",
7097 => "0000000000000000",7098 => "0000000000000000",
7099 => "0000000000000000",7100 => "0000000000000000",
7101 => "0000000000000000",7102 => "0000000000000000",
7103 => "0000000000000000",7104 => "0000000000000000",
7105 => "0000000000000000",7106 => "0000000000000000",
7107 => "0000000000000000",7108 => "0000000000000000",
7109 => "0000000000000000",7110 => "0000000000000000",
7111 => "0000000000000000",7112 => "0000000000000000",
7113 => "0000000000000000",7114 => "0000000000000000",
7115 => "0000000000000000",7116 => "0000000000000000",
7117 => "0000000000000000",7118 => "0000000000000000",
7119 => "0000000000000000",7120 => "0000000000000000",
7121 => "0000000000000000",7122 => "0000000000000000",
7123 => "0000000000000000",7124 => "0000000000000000",
7125 => "0000000000000000",7126 => "0000000000000000",
7127 => "0000000000000000",7128 => "0000000000000000",
7129 => "0000000000000000",7130 => "0000000000000000",
7131 => "0000000000000000",7132 => "0000000000000000",
7133 => "0000000000000000",7134 => "0000000000000000",
7135 => "0000000000000000",7136 => "0000000000000000",
7137 => "0000000000000000",7138 => "0000000000000000",
7139 => "0000000000000000",7140 => "0000000000000000",
7141 => "0000000000000000",7142 => "0000000000000000",
7143 => "0000000000000000",7144 => "0000000000000000",
7145 => "0000000000000000",7146 => "0000000000000000",
7147 => "0000000000000000",7148 => "0000000000000000",
7149 => "0000000000000000",7150 => "0000000000000000",
7151 => "0000000000000000",7152 => "0000000000000000",
7153 => "0000000000000000",7154 => "0000000000000000",
7155 => "0000000000000000",7156 => "0000000000000000",
7157 => "0000000000000000",7158 => "0000000000000000",
7159 => "0000000000000000",7160 => "0000000000000000",
7161 => "0000000000000000",7162 => "0000000000000000",
7163 => "0000000000000000",7164 => "0000000000000000",
7165 => "0000000000000000",7166 => "0000000000000000",
7167 => "0000000000000000",7168 => "0000000000000000",
7169 => "0000000000000000",7170 => "0000000000000000",
7171 => "0000000000000000",7172 => "0000000000000000",
7173 => "0000000000000000",7174 => "0000000000000000",
7175 => "0000000000000000",7176 => "0000000000000000",
7177 => "0000000000000000",7178 => "0000000000000000",
7179 => "0000000000000000",7180 => "0000000000000000",
7181 => "0000000000000000",7182 => "0000000000000000",
7183 => "0000000000000000",7184 => "0000000000000000",
7185 => "0000000000000000",7186 => "0000000000000000",
7187 => "0000000000000000",7188 => "0000000000000000",
7189 => "0000000000000000",7190 => "0000000000000000",
7191 => "0000000000000000",7192 => "0000000000000000",
7193 => "0000000000000000",7194 => "0000000000000000",
7195 => "0000000000000000",7196 => "0000000000000000",
7197 => "0000000000000000",7198 => "0000000000000000",
7199 => "0000000000000000",7200 => "0000000000000000",
7201 => "0000000000000000",7202 => "0000000000000000",
7203 => "0000000000000000",7204 => "0000000000000000",
7205 => "0000000000000000",7206 => "0000000000000000",
7207 => "0000000000000000",7208 => "0000000000000000",
7209 => "0000000000000000",7210 => "0000000000000000",
7211 => "0000000000000000",7212 => "0000000000000000",
7213 => "0000000000000000",7214 => "0000000000000000",
7215 => "0000000000000000",7216 => "0000000000000000",
7217 => "0000000000000000",7218 => "0000000000000000",
7219 => "0000000000000000",7220 => "0000000000000000",
7221 => "0000000000000000",7222 => "0000000000000000",
7223 => "0000000000000000",7224 => "0000000000000000",
7225 => "0000000000000000",7226 => "0000000000000000",
7227 => "0000000000000000",7228 => "0000000000000000",
7229 => "0000000000000000",7230 => "0000000000000000",
7231 => "0000000000000000",7232 => "0000000000000000",
7233 => "0000000000000000",7234 => "0000000000000000",
7235 => "0000000000000000",7236 => "0000000000000000",
7237 => "0000000000000000",7238 => "0000000000000000",
7239 => "0000000000000000",7240 => "0000000000000000",
7241 => "0000000000000000",7242 => "0000000000000000",
7243 => "0000000000000000",7244 => "0000000000000000",
7245 => "0000000000000000",7246 => "0000000000000000",
7247 => "0000000000000000",7248 => "0000000000000000",
7249 => "0000000000000000",7250 => "0000000000000000",
7251 => "0000000000000000",7252 => "0000000000000000",
7253 => "0000000000000000",7254 => "0000000000000000",
7255 => "0000000000000000",7256 => "0000000000000000",
7257 => "0000000000000000",7258 => "0000000000000000",
7259 => "0000000000000000",7260 => "0000000000000000",
7261 => "0000000000000000",7262 => "0000000000000000",
7263 => "0000000000000000",7264 => "0000000000000000",
7265 => "0000000000000000",7266 => "0000000000000000",
7267 => "0000000000000000",7268 => "0000000000000000",
7269 => "0000000000000000",7270 => "0000000000000000",
7271 => "0000000000000000",7272 => "0000000000000000",
7273 => "0000000000000000",7274 => "0000000000000000",
7275 => "0000000000000000",7276 => "0000000000000000",
7277 => "0000000000000000",7278 => "0000000000000000",
7279 => "0000000000000000",7280 => "0000000000000000",
7281 => "0000000000000000",7282 => "0000000000000000",
7283 => "0000000000000000",7284 => "0000000000000000",
7285 => "0000000000000000",7286 => "0000000000000000",
7287 => "0000000000000000",7288 => "0000000000000000",
7289 => "0000000000000000",7290 => "0000000000000000",
7291 => "0000000000000000",7292 => "0000000000000000",
7293 => "0000000000000000",7294 => "0000000000000000",
7295 => "0000000000000000",7296 => "0000000000000000",
7297 => "0000000000000000",7298 => "0000000000000000",
7299 => "0000000000000000",7300 => "0000000000000000",
7301 => "0000000000000000",7302 => "0000000000000000",
7303 => "0000000000000000",7304 => "0000000000000000",
7305 => "0000000000000000",7306 => "0000000000000000",
7307 => "0000000000000000",7308 => "0000000000000000",
7309 => "0000000000000000",7310 => "0000000000000000",
7311 => "0000000000000000",7312 => "0000000000000000",
7313 => "0000000000000000",7314 => "0000000000000000",
7315 => "0000000000000000",7316 => "0000000000000000",
7317 => "0000000000000000",7318 => "0000000000000000",
7319 => "0000000000000000",7320 => "0000000000000000",
7321 => "0000000000000000",7322 => "0000000000000000",
7323 => "0000000000000000",7324 => "0000000000000000",
7325 => "0000000000000000",7326 => "0000000000000000",
7327 => "0000000000000000",7328 => "0000000000000000",
7329 => "0000000000000000",7330 => "0000000000000000",
7331 => "0000000000000000",7332 => "0000000000000000",
7333 => "0000000000000000",7334 => "0000000000000000",
7335 => "0000000000000000",7336 => "0000000000000000",
7337 => "0000000000000000",7338 => "0000000000000000",
7339 => "0000000000000000",7340 => "0000000000000000",
7341 => "0000000000000000",7342 => "0000000000000000",
7343 => "0000000000000000",7344 => "0000000000000000",
7345 => "0000000000000000",7346 => "0000000000000000",
7347 => "0000000000000000",7348 => "0000000000000000",
7349 => "0000000000000000",7350 => "0000000000000000",
7351 => "0000000000000000",7352 => "0000000000000000",
7353 => "0000000000000000",7354 => "0000000000000000",
7355 => "0000000000000000",7356 => "0000000000000000",
7357 => "0000000000000000",7358 => "0000000000000000",
7359 => "0000000000000000",7360 => "0000000000000000",
7361 => "0000000000000000",7362 => "0000000000000000",
7363 => "0000000000000000",7364 => "0000000000000000",
7365 => "0000000000000000",7366 => "0000000000000000",
7367 => "0000000000000000",7368 => "0000000000000000",
7369 => "0000000000000000",7370 => "0000000000000000",
7371 => "0000000000000000",7372 => "0000000000000000",
7373 => "0000000000000000",7374 => "0000000000000000",
7375 => "0000000000000000",7376 => "0000000000000000",
7377 => "0000000000000000",7378 => "0000000000000000",
7379 => "0000000000000000",7380 => "0000000000000000",
7381 => "0000000000000000",7382 => "0000000000000000",
7383 => "0000000000000000",7384 => "0000000000000000",
7385 => "0000000000000000",7386 => "0000000000000000",
7387 => "0000000000000000",7388 => "0000000000000000",
7389 => "0000000000000000",7390 => "0000000000000000",
7391 => "0000000000000000",7392 => "0000000000000000",
7393 => "0000000000000000",7394 => "0000000000000000",
7395 => "0000000000000000",7396 => "0000000000000000",
7397 => "0000000000000000",7398 => "0000000000000000",
7399 => "0000000000000000",7400 => "0000000000000000",
7401 => "0000000000000000",7402 => "0000000000000000",
7403 => "0000000000000000",7404 => "0000000000000000",
7405 => "0000000000000000",7406 => "0000000000000000",
7407 => "0000000000000000",7408 => "0000000000000000",
7409 => "0000000000000000",7410 => "0000000000000000",
7411 => "0000000000000000",7412 => "0000000000000000",
7413 => "0000000000000000",7414 => "0000000000000000",
7415 => "0000000000000000",7416 => "0000000000000000",
7417 => "0000000000000000",7418 => "0000000000000000",
7419 => "0000000000000000",7420 => "0000000000000000",
7421 => "0000000000000000",7422 => "0000000000000000",
7423 => "0000000000000000",7424 => "0000000000000000",
7425 => "0000000000000000",7426 => "0000000000000000",
7427 => "0000000000000000",7428 => "0000000000000000",
7429 => "0000000000000000",7430 => "0000000000000000",
7431 => "0000000000000000",7432 => "0000000000000000",
7433 => "0000000000000000",7434 => "0000000000000000",
7435 => "0000000000000000",7436 => "0000000000000000",
7437 => "0000000000000000",7438 => "0000000000000000",
7439 => "0000000000000000",7440 => "0000000000000000",
7441 => "0000000000000000",7442 => "0000000000000000",
7443 => "0000000000000000",7444 => "0000000000000000",
7445 => "0000000000000000",7446 => "0000000000000000",
7447 => "0000000000000000",7448 => "0000000000000000",
7449 => "0000000000000000",7450 => "0000000000000000",
7451 => "0000000000000000",7452 => "0000000000000000",
7453 => "0000000000000000",7454 => "0000000000000000",
7455 => "0000000000000000",7456 => "0000000000000000",
7457 => "0000000000000000",7458 => "0000000000000000",
7459 => "0000000000000000",7460 => "0000000000000000",
7461 => "0000000000000000",7462 => "0000000000000000",
7463 => "0000000000000000",7464 => "0000000000000000",
7465 => "0000000000000000",7466 => "0000000000000000",
7467 => "0000000000000000",7468 => "0000000000000000",
7469 => "0000000000000000",7470 => "0000000000000000",
7471 => "0000000000000000",7472 => "0000000000000000",
7473 => "0000000000000000",7474 => "0000000000000000",
7475 => "0000000000000000",7476 => "0000000000000000",
7477 => "0000000000000000",7478 => "0000000000000000",
7479 => "0000000000000000",7480 => "0000000000000000",
7481 => "0000000000000000",7482 => "0000000000000000",
7483 => "0000000000000000",7484 => "0000000000000000",
7485 => "0000000000000000",7486 => "0000000000000000",
7487 => "0000000000000000",7488 => "0000000000000000",
7489 => "0000000000000000",7490 => "0000000000000000",
7491 => "0000000000000000",7492 => "0000000000000000",
7493 => "0000000000000000",7494 => "0000000000000000",
7495 => "0000000000000000",7496 => "0000000000000000",
7497 => "0000000000000000",7498 => "0000000000000000",
7499 => "0000000000000000",7500 => "0000000000000000",
7501 => "0000000000000000",7502 => "0000000000000000",
7503 => "0000000000000000",7504 => "0000000000000000",
7505 => "0000000000000000",7506 => "0000000000000000",
7507 => "0000000000000000",7508 => "0000000000000000",
7509 => "0000000000000000",7510 => "0000000000000000",
7511 => "0000000000000000",7512 => "0000000000000000",
7513 => "0000000000000000",7514 => "0000000000000000",
7515 => "0000000000000000",7516 => "0000000000000000",
7517 => "0000000000000000",7518 => "0000000000000000",
7519 => "0000000000000000",7520 => "0000000000000000",
7521 => "0000000000000000",7522 => "0000000000000000",
7523 => "0000000000000000",7524 => "0000000000000000",
7525 => "0000000000000000",7526 => "0000000000000000",
7527 => "0000000000000000",7528 => "0000000000000000",
7529 => "0000000000000000",7530 => "0000000000000000",
7531 => "0000000000000000",7532 => "0000000000000000",
7533 => "0000000000000000",7534 => "0000000000000000",
7535 => "0000000000000000",7536 => "0000000000000000",
7537 => "0000000000000000",7538 => "0000000000000000",
7539 => "0000000000000000",7540 => "0000000000000000",
7541 => "0000000000000000",7542 => "0000000000000000",
7543 => "0000000000000000",7544 => "0000000000000000",
7545 => "0000000000000000",7546 => "0000000000000000",
7547 => "0000000000000000",7548 => "0000000000000000",
7549 => "0000000000000000",7550 => "0000000000000000",
7551 => "0000000000000000",7552 => "0000000000000000",
7553 => "0000000000000000",7554 => "0000000000000000",
7555 => "0000000000000000",7556 => "0000000000000000",
7557 => "0000000000000000",7558 => "0000000000000000",
7559 => "0000000000000000",7560 => "0000000000000000",
7561 => "0000000000000000",7562 => "0000000000000000",
7563 => "0000000000000000",7564 => "0000000000000000",
7565 => "0000000000000000",7566 => "0000000000000000",
7567 => "0000000000000000",7568 => "0000000000000000",
7569 => "0000000000000000",7570 => "0000000000000000",
7571 => "0000000000000000",7572 => "0000000000000000",
7573 => "0000000000000000",7574 => "0000000000000000",
7575 => "0000000000000000",7576 => "0000000000000000",
7577 => "0000000000000000",7578 => "0000000000000000",
7579 => "0000000000000000",7580 => "0000000000000000",
7581 => "0000000000000000",7582 => "0000000000000000",
7583 => "0000000000000000",7584 => "0000000000000000",
7585 => "0000000000000000",7586 => "0000000000000000",
7587 => "0000000000000000",7588 => "0000000000000000",
7589 => "0000000000000000",7590 => "0000000000000000",
7591 => "0000000000000000",7592 => "0000000000000000",
7593 => "0000000000000000",7594 => "0000000000000000",
7595 => "0000000000000000",7596 => "0000000000000000",
7597 => "0000000000000000",7598 => "0000000000000000",
7599 => "0000000000000000",7600 => "0000000000000000",
7601 => "0000000000000000",7602 => "0000000000000000",
7603 => "0000000000000000",7604 => "0000000000000000",
7605 => "0000000000000000",7606 => "0000000000000000",
7607 => "0000000000000000",7608 => "0000000000000000",
7609 => "0000000000000000",7610 => "0000000000000000",
7611 => "0000000000000000",7612 => "0000000000000000",
7613 => "0000000000000000",7614 => "0000000000000000",
7615 => "0000000000000000",7616 => "0000000000000000",
7617 => "0000000000000000",7618 => "0000000000000000",
7619 => "0000000000000000",7620 => "0000000000000000",
7621 => "0000000000000000",7622 => "0000000000000000",
7623 => "0000000000000000",7624 => "0000000000000000",
7625 => "0000000000000000",7626 => "0000000000000000",
7627 => "0000000000000000",7628 => "0000000000000000",
7629 => "0000000000000000",7630 => "0000000000000000",
7631 => "0000000000000000",7632 => "0000000000000000",
7633 => "0000000000000000",7634 => "0000000000000000",
7635 => "0000000000000000",7636 => "0000000000000000",
7637 => "0000000000000000",7638 => "0000000000000000",
7639 => "0000000000000000",7640 => "0000000000000000",
7641 => "0000000000000000",7642 => "0000000000000000",
7643 => "0000000000000000",7644 => "0000000000000000",
7645 => "0000000000000000",7646 => "0000000000000000",
7647 => "0000000000000000",7648 => "0000000000000000",
7649 => "0000000000000000",7650 => "0000000000000000",
7651 => "0000000000000000",7652 => "0000000000000000",
7653 => "0000000000000000",7654 => "0000000000000000",
7655 => "0000000000000000",7656 => "0000000000000000",
7657 => "0000000000000000",7658 => "0000000000000000",
7659 => "0000000000000000",7660 => "0000000000000000",
7661 => "0000000000000000",7662 => "0000000000000000",
7663 => "0000000000000000",7664 => "0000000000000000",
7665 => "0000000000000000",7666 => "0000000000000000",
7667 => "0000000000000000",7668 => "0000000000000000",
7669 => "0000000000000000",7670 => "0000000000000000",
7671 => "0000000000000000",7672 => "0000000000000000",
7673 => "0000000000000000",7674 => "0000000000000000",
7675 => "0000000000000000",7676 => "0000000000000000",
7677 => "0000000000000000",7678 => "0000000000000000",
7679 => "0000000000000000",7680 => "0000000000000000",
7681 => "0000000000000000",7682 => "0000000000000000",
7683 => "0000000000000000",7684 => "0000000000000000",
7685 => "0000000000000000",7686 => "0000000000000000",
7687 => "0000000000000000",7688 => "0000000000000000",
7689 => "0000000000000000",7690 => "0000000000000000",
7691 => "0000000000000000",7692 => "0000000000000000",
7693 => "0000000000000000",7694 => "0000000000000000",
7695 => "0000000000000000",7696 => "0000000000000000",
7697 => "0000000000000000",7698 => "0000000000000000",
7699 => "0000000000000000",7700 => "0000000000000000",
7701 => "0000000000000000",7702 => "0000000000000000",
7703 => "0000000000000000",7704 => "0000000000000000",
7705 => "0000000000000000",7706 => "0000000000000000",
7707 => "0000000000000000",7708 => "0000000000000000",
7709 => "0000000000000000",7710 => "0000000000000000",
7711 => "0000000000000000",7712 => "0000000000000000",
7713 => "0000000000000000",7714 => "0000000000000000",
7715 => "0000000000000000",7716 => "0000000000000000",
7717 => "0000000000000000",7718 => "0000000000000000",
7719 => "0000000000000000",7720 => "0000000000000000",
7721 => "0000000000000000",7722 => "0000000000000000",
7723 => "0000000000000000",7724 => "0000000000000000",
7725 => "0000000000000000",7726 => "0000000000000000",
7727 => "0000000000000000",7728 => "0000000000000000",
7729 => "0000000000000000",7730 => "0000000000000000",
7731 => "0000000000000000",7732 => "0000000000000000",
7733 => "0000000000000000",7734 => "0000000000000000",
7735 => "0000000000000000",7736 => "0000000000000000",
7737 => "0000000000000000",7738 => "0000000000000000",
7739 => "0000000000000000",7740 => "0000000000000000",
7741 => "0000000000000000",7742 => "0000000000000000",
7743 => "0000000000000000",7744 => "0000000000000000",
7745 => "0000000000000000",7746 => "0000000000000000",
7747 => "0000000000000000",7748 => "0000000000000000",
7749 => "0000000000000000",7750 => "0000000000000000",
7751 => "0000000000000000",7752 => "0000000000000000",
7753 => "0000000000000000",7754 => "0000000000000000",
7755 => "0000000000000000",7756 => "0000000000000000",
7757 => "0000000000000000",7758 => "0000000000000000",
7759 => "0000000000000000",7760 => "0000000000000000",
7761 => "0000000000000000",7762 => "0000000000000000",
7763 => "0000000000000000",7764 => "0000000000000000",
7765 => "0000000000000000",7766 => "0000000000000000",
7767 => "0000000000000000",7768 => "0000000000000000",
7769 => "0000000000000000",7770 => "0000000000000000",
7771 => "0000000000000000",7772 => "0000000000000000",
7773 => "0000000000000000",7774 => "0000000000000000",
7775 => "0000000000000000",7776 => "0000000000000000",
7777 => "0000000000000000",7778 => "0000000000000000",
7779 => "0000000000000000",7780 => "0000000000000000",
7781 => "0000000000000000",7782 => "0000000000000000",
7783 => "0000000000000000",7784 => "0000000000000000",
7785 => "0000000000000000",7786 => "0000000000000000",
7787 => "0000000000000000",7788 => "0000000000000000",
7789 => "0000000000000000",7790 => "0000000000000000",
7791 => "0000000000000000",7792 => "0000000000000000",
7793 => "0000000000000000",7794 => "0000000000000000",
7795 => "0000000000000000",7796 => "0000000000000000",
7797 => "0000000000000000",7798 => "0000000000000000",
7799 => "0000000000000000",7800 => "0000000000000000",
7801 => "0000000000000000",7802 => "0000000000000000",
7803 => "0000000000000000",7804 => "0000000000000000",
7805 => "0000000000000000",7806 => "0000000000000000",
7807 => "0000000000000000",7808 => "0000000000000000",
7809 => "0000000000000000",7810 => "0000000000000000",
7811 => "0000000000000000",7812 => "0000000000000000",
7813 => "0000000000000000",7814 => "0000000000000000",
7815 => "0000000000000000",7816 => "0000000000000000",
7817 => "0000000000000000",7818 => "0000000000000000",
7819 => "0000000000000000",7820 => "0000000000000000",
7821 => "0000000000000000",7822 => "0000000000000000",
7823 => "0000000000000000",7824 => "0000000000000000",
7825 => "0000000000000000",7826 => "0000000000000000",
7827 => "0000000000000000",7828 => "0000000000000000",
7829 => "0000000000000000",7830 => "0000000000000000",
7831 => "0000000000000000",7832 => "0000000000000000",
7833 => "0000000000000000",7834 => "0000000000000000",
7835 => "0000000000000000",7836 => "0000000000000000",
7837 => "0000000000000000",7838 => "0000000000000000",
7839 => "0000000000000000",7840 => "0000000000000000",
7841 => "0000000000000000",7842 => "0000000000000000",
7843 => "0000000000000000",7844 => "0000000000000000",
7845 => "0000000000000000",7846 => "0000000000000000",
7847 => "0000000000000000",7848 => "0000000000000000",
7849 => "0000000000000000",7850 => "0000000000000000",
7851 => "0000000000000000",7852 => "0000000000000000",
7853 => "0000000000000000",7854 => "0000000000000000",
7855 => "0000000000000000",7856 => "0000000000000000",
7857 => "0000000000000000",7858 => "0000000000000000",
7859 => "0000000000000000",7860 => "0000000000000000",
7861 => "0000000000000000",7862 => "0000000000000000",
7863 => "0000000000000000",7864 => "0000000000000000",
7865 => "0000000000000000",7866 => "0000000000000000",
7867 => "0000000000000000",7868 => "0000000000000000",
7869 => "0000000000000000",7870 => "0000000000000000",
7871 => "0000000000000000",7872 => "0000000000000000",
7873 => "0000000000000000",7874 => "0000000000000000",
7875 => "0000000000000000",7876 => "0000000000000000",
7877 => "0000000000000000",7878 => "0000000000000000",
7879 => "0000000000000000",7880 => "0000000000000000",
7881 => "0000000000000000",7882 => "0000000000000000",
7883 => "0000000000000000",7884 => "0000000000000000",
7885 => "0000000000000000",7886 => "0000000000000000",
7887 => "0000000000000000",7888 => "0000000000000000",
7889 => "0000000000000000",7890 => "0000000000000000",
7891 => "0000000000000000",7892 => "0000000000000000",
7893 => "0000000000000000",7894 => "0000000000000000",
7895 => "0000000000000000",7896 => "0000000000000000",
7897 => "0000000000000000",7898 => "0000000000000000",
7899 => "0000000000000000",7900 => "0000000000000000",
7901 => "0000000000000000",7902 => "0000000000000000",
7903 => "0000000000000000",7904 => "0000000000000000",
7905 => "0000000000000000",7906 => "0000000000000000",
7907 => "0000000000000000",7908 => "0000000000000000",
7909 => "0000000000000000",7910 => "0000000000000000",
7911 => "0000000000000000",7912 => "0000000000000000",
7913 => "0000000000000000",7914 => "0000000000000000",
7915 => "0000000000000000",7916 => "0000000000000000",
7917 => "0000000000000000",7918 => "0000000000000000",
7919 => "0000000000000000",7920 => "0000000000000000",
7921 => "0000000000000000",7922 => "0000000000000000",
7923 => "0000000000000000",7924 => "0000000000000000",
7925 => "0000000000000000",7926 => "0000000000000000",
7927 => "0000000000000000",7928 => "0000000000000000",
7929 => "0000000000000000",7930 => "0000000000000000",
7931 => "0000000000000000",7932 => "0000000000000000",
7933 => "0000000000000000",7934 => "0000000000000000",
7935 => "0000000000000000",7936 => "0000000000000000",
7937 => "0000000000000000",7938 => "0000000000000000",
7939 => "0000000000000000",7940 => "0000000000000000",
7941 => "0000000000000000",7942 => "0000000000000000",
7943 => "0000000000000000",7944 => "0000000000000000",
7945 => "0000000000000000",7946 => "0000000000000000",
7947 => "0000000000000000",7948 => "0000000000000000",
7949 => "0000000000000000",7950 => "0000000000000000",
7951 => "0000000000000000",7952 => "0000000000000000",
7953 => "0000000000000000",7954 => "0000000000000000",
7955 => "0000000000000000",7956 => "0000000000000000",
7957 => "0000000000000000",7958 => "0000000000000000",
7959 => "0000000000000000",7960 => "0000000000000000",
7961 => "0000000000000000",7962 => "0000000000000000",
7963 => "0000000000000000",7964 => "0000000000000000",
7965 => "0000000000000000",7966 => "0000000000000000",
7967 => "0000000000000000",7968 => "0000000000000000",
7969 => "0000000000000000",7970 => "0000000000000000",
7971 => "0000000000000000",7972 => "0000000000000000",
7973 => "0000000000000000",7974 => "0000000000000000",
7975 => "0000000000000000",7976 => "0000000000000000",
7977 => "0000000000000000",7978 => "0000000000000000",
7979 => "0000000000000000",7980 => "0000000000000000",
7981 => "0000000000000000",7982 => "0000000000000000",
7983 => "0000000000000000",7984 => "0000000000000000",
7985 => "0000000000000000",7986 => "0000000000000000",
7987 => "0000000000000000",7988 => "0000000000000000",
7989 => "0000000000000000",7990 => "0000000000000000",
7991 => "0000000000000000",7992 => "0000000000000000",
7993 => "0000000000000000",7994 => "0000000000000000",
7995 => "0000000000000000",7996 => "0000000000000000",
7997 => "0000000000000000",7998 => "0000000000000000",
7999 => "0000000000000000",8000 => "0000000000000000",
8001 => "0000000000000000",8002 => "0000000000000000",
8003 => "0000000000000000",8004 => "0000000000000000",
8005 => "0000000000000000",8006 => "0000000000000000",
8007 => "0000000000000000",8008 => "0000000000000000",
8009 => "0000000000000000",8010 => "0000000000000000",
8011 => "0000000000000000",8012 => "0000000000000000",
8013 => "0000000000000000",8014 => "0000000000000000",
8015 => "0000000000000000",8016 => "0000000000000000",
8017 => "0000000000000000",8018 => "0000000000000000",
8019 => "0000000000000000",8020 => "0000000000000000",
8021 => "0000000000000000",8022 => "0000000000000000",
8023 => "0000000000000000",8024 => "0000000000000000",
8025 => "0000000000000000",8026 => "0000000000000000",
8027 => "0000000000000000",8028 => "0000000000000000",
8029 => "0000000000000000",8030 => "0000000000000000",
8031 => "0000000000000000",8032 => "0000000000000000",
8033 => "0000000000000000",8034 => "0000000000000000",
8035 => "0000000000000000",8036 => "0000000000000000",
8037 => "0000000000000000",8038 => "0000000000000000",
8039 => "0000000000000000",8040 => "0000000000000000",
8041 => "0000000000000000",8042 => "0000000000000000",
8043 => "0000000000000000",8044 => "0000000000000000",
8045 => "0000000000000000",8046 => "0000000000000000",
8047 => "0000000000000000",8048 => "0000000000000000",
8049 => "0000000000000000",8050 => "0000000000000000",
8051 => "0000000000000000",8052 => "0000000000000000",
8053 => "0000000000000000",8054 => "0000000000000000",
8055 => "0000000000000000",8056 => "0000000000000000",
8057 => "0000000000000000",8058 => "0000000000000000",
8059 => "0000000000000000",8060 => "0000000000000000",
8061 => "0000000000000000",8062 => "0000000000000000",
8063 => "0000000000000000",8064 => "0000000000000000",
8065 => "0000000000000000",8066 => "0000000000000000",
8067 => "0000000000000000",8068 => "0000000000000000",
8069 => "0000000000000000",8070 => "0000000000000000",
8071 => "0000000000000000",8072 => "0000000000000000",
8073 => "0000000000000000",8074 => "0000000000000000",
8075 => "0000000000000000",8076 => "0000000000000000",
8077 => "0000000000000000",8078 => "0000000000000000",
8079 => "0000000000000000",8080 => "0000000000000000",
8081 => "0000000000000000",8082 => "0000000000000000",
8083 => "0000000000000000",8084 => "0000000000000000",
8085 => "0000000000000000",8086 => "0000000000000000",
8087 => "0000000000000000",8088 => "0000000000000000",
8089 => "0000000000000000",8090 => "0000000000000000",
8091 => "0000000000000000",8092 => "0000000000000000",
8093 => "0000000000000000",8094 => "0000000000000000",
8095 => "0000000000000000",8096 => "0000000000000000",
8097 => "0000000000000000",8098 => "0000000000000000",
8099 => "0000000000000000",8100 => "0000000000000000",
8101 => "0000000000000000",8102 => "0000000000000000",
8103 => "0000000000000000",8104 => "0000000000000000",
8105 => "0000000000000000",8106 => "0000000000000000",
8107 => "0000000000000000",8108 => "0000000000000000",
8109 => "0000000000000000",8110 => "0000000000000000",
8111 => "0000000000000000",8112 => "0000000000000000",
8113 => "0000000000000000",8114 => "0000000000000000",
8115 => "0000000000000000",8116 => "0000000000000000",
8117 => "0000000000000000",8118 => "0000000000000000",
8119 => "0000000000000000",8120 => "0000000000000000",
8121 => "0000000000000000",8122 => "0000000000000000",
8123 => "0000000000000000",8124 => "0000000000000000",
8125 => "0000000000000000",8126 => "0000000000000000",
8127 => "0000000000000000",8128 => "0000000000000000",
8129 => "0000000000000000",8130 => "0000000000000000",
8131 => "0000000000000000",8132 => "0000000000000000",
8133 => "0000000000000000",8134 => "0000000000000000",
8135 => "0000000000000000",8136 => "0000000000000000",
8137 => "0000000000000000",8138 => "0000000000000000",
8139 => "0000000000000000",8140 => "0000000000000000",
8141 => "0000000000000000",8142 => "0000000000000000",
8143 => "0000000000000000",8144 => "0000000000000000",
8145 => "0000000000000000",8146 => "0000000000000000",
8147 => "0000000000000000",8148 => "0000000000000000",
8149 => "0000000000000000",8150 => "0000000000000000",
8151 => "0000000000000000",8152 => "0000000000000000",
8153 => "0000000000000000",8154 => "0000000000000000",
8155 => "0000000000000000",8156 => "0000000000000000",
8157 => "0000000000000000",8158 => "0000000000000000",
8159 => "0000000000000000",8160 => "0000000000000000",
8161 => "0000000000000000",8162 => "0000000000000000",
8163 => "0000000000000000",8164 => "0000000000000000",
8165 => "0000000000000000",8166 => "0000000000000000",
8167 => "0000000000000000",8168 => "0000000000000000",
8169 => "0000000000000000",8170 => "0000000000000000",
8171 => "0000000000000000",8172 => "0000000000000000",
8173 => "0000000000000000",8174 => "0000000000000000",
8175 => "0000000000000000",8176 => "0000000000000000",
8177 => "0000000000000000",8178 => "0000000000000000",
8179 => "0000000000000000",8180 => "0000000000000000",
8181 => "0000000000000000",8182 => "0000000000000000",
8183 => "0000000000000000",8184 => "0000000000000000",
8185 => "0000000000000000",8186 => "0000000000000000",
8187 => "0000000000000000",8188 => "0000000000000000",
8189 => "0000000000000000",8190 => "0000000000000000",
8191 => "0000000000000000",8192 => "0000000000000000",
8193 => "0000000000000000",8194 => "0000000000000000",
8195 => "0000000000000000",8196 => "0000000000000000",
8197 => "0000000000000000",8198 => "0000000000000000",
8199 => "0000000000000000",8200 => "0000000000000000",
8201 => "0000000000000000",8202 => "0000000000000000",
8203 => "0000000000000000",8204 => "0000000000000000",
8205 => "0000000000000000",8206 => "0000000000000000",
8207 => "0000000000000000",8208 => "0000000000000000",
8209 => "0000000000000000",8210 => "0000000000000000",
8211 => "0000000000000000",8212 => "0000000000000000",
8213 => "0000000000000000",8214 => "0000000000000000",
8215 => "0000000000000000",8216 => "0000000000000000",
8217 => "0000000000000000",8218 => "0000000000000000",
8219 => "0000000000000000",8220 => "0000000000000000",
8221 => "0000000000000000",8222 => "0000000000000000",
8223 => "0000000000000000",8224 => "0000000000000000",
8225 => "0000000000000000",8226 => "0000000000000000",
8227 => "0000000000000000",8228 => "0000000000000000",
8229 => "0000000000000000",8230 => "0000000000000000",
8231 => "0000000000000000",8232 => "0000000000000000",
8233 => "0000000000000000",8234 => "0000000000000000",
8235 => "0000000000000000",8236 => "0000000000000000",
8237 => "0000000000000000",8238 => "0000000000000000",
8239 => "0000000000000000",8240 => "0000000000000000",
8241 => "0000000000000000",8242 => "0000000000000000",
8243 => "0000000000000000",8244 => "0000000000000000",
8245 => "0000000000000000",8246 => "0000000000000000",
8247 => "0000000000000000",8248 => "0000000000000000",
8249 => "0000000000000000",8250 => "0000000000000000",
8251 => "0000000000000000",8252 => "0000000000000000",
8253 => "0000000000000000",8254 => "0000000000000000",
8255 => "0000000000000000",8256 => "0000000000000000",
8257 => "0000000000000000",8258 => "0000000000000000",
8259 => "0000000000000000",8260 => "0000000000000000",
8261 => "0000000000000000",8262 => "0000000000000000",
8263 => "0000000000000000",8264 => "0000000000000000",
8265 => "0000000000000000",8266 => "0000000000000000",
8267 => "0000000000000000",8268 => "0000000000000000",
8269 => "0000000000000000",8270 => "0000000000000000",
8271 => "0000000000000000",8272 => "0000000000000000",
8273 => "0000000000000000",8274 => "0000000000000000",
8275 => "0000000000000000",8276 => "0000000000000000",
8277 => "0000000000000000",8278 => "0000000000000000",
8279 => "0000000000000000",8280 => "0000000000000000",
8281 => "0000000000000000",8282 => "0000000000000000",
8283 => "0000000000000000",8284 => "0000000000000000",
8285 => "0000000000000000",8286 => "0000000000000000",
8287 => "0000000000000000",8288 => "0000000000000000",
8289 => "0000000000000000",8290 => "0000000000000000",
8291 => "0000000000000000",8292 => "0000000000000000",
8293 => "0000000000000000",8294 => "0000000000000000",
8295 => "0000000000000000",8296 => "0000000000000000",
8297 => "0000000000000000",8298 => "0000000000000000",
8299 => "0000000000000000",8300 => "0000000000000000",
8301 => "0000000000000000",8302 => "0000000000000000",
8303 => "0000000000000000",8304 => "0000000000000000",
8305 => "0000000000000000",8306 => "0000000000000000",
8307 => "0000000000000000",8308 => "0000000000000000",
8309 => "0000000000000000",8310 => "0000000000000000",
8311 => "0000000000000000",8312 => "0000000000000000",
8313 => "0000000000000000",8314 => "0000000000000000",
8315 => "0000000000000000",8316 => "0000000000000000",
8317 => "0000000000000000",8318 => "0000000000000000",
8319 => "0000000000000000",8320 => "0000000000000000",
8321 => "0000000000000000",8322 => "0000000000000000",
8323 => "0000000000000000",8324 => "0000000000000000",
8325 => "0000000000000000",8326 => "0000000000000000",
8327 => "0000000000000000",8328 => "0000000000000000",
8329 => "0000000000000000",8330 => "0000000000000000",
8331 => "0000000000000000",8332 => "0000000000000000",
8333 => "0000000000000000",8334 => "0000000000000000",
8335 => "0000000000000000",8336 => "0000000000000000",
8337 => "0000000000000000",8338 => "0000000000000000",
8339 => "0000000000000000",8340 => "0000000000000000",
8341 => "0000000000000000",8342 => "0000000000000000",
8343 => "0000000000000000",8344 => "0000000000000000",
8345 => "0000000000000000",8346 => "0000000000000000",
8347 => "0000000000000000",8348 => "0000000000000000",
8349 => "0000000000000000",8350 => "0000000000000000",
8351 => "0000000000000000",8352 => "0000000000000000",
8353 => "0000000000000000",8354 => "0000000000000000",
8355 => "0000000000000000",8356 => "0000000000000000",
8357 => "0000000000000000",8358 => "0000000000000000",
8359 => "0000000000000000",8360 => "0000000000000000",
8361 => "0000000000000000",8362 => "0000000000000000",
8363 => "0000000000000000",8364 => "0000000000000000",
8365 => "0000000000000000",8366 => "0000000000000000",
8367 => "0000000000000000",8368 => "0000000000000000",
8369 => "0000000000000000",8370 => "0000000000000000",
8371 => "0000000000000000",8372 => "0000000000000000",
8373 => "0000000000000000",8374 => "0000000000000000",
8375 => "0000000000000000",8376 => "0000000000000000",
8377 => "0000000000000000",8378 => "0000000000000000",
8379 => "0000000000000000",8380 => "0000000000000000",
8381 => "0000000000000000",8382 => "0000000000000000",
8383 => "0000000000000000",8384 => "0000000000000000",
8385 => "0000000000000000",8386 => "0000000000000000",
8387 => "0000000000000000",8388 => "0000000000000000",
8389 => "0000000000000000",8390 => "0000000000000000",
8391 => "0000000000000000",8392 => "0000000000000000",
8393 => "0000000000000000",8394 => "0000000000000000",
8395 => "0000000000000000",8396 => "0000000000000000",
8397 => "0000000000000000",8398 => "0000000000000000",
8399 => "0000000000000000",8400 => "0000000000000000",
8401 => "0000000000000000",8402 => "0000000000000000",
8403 => "0000000000000000",8404 => "0000000000000000",
8405 => "0000000000000000",8406 => "0000000000000000",
8407 => "0000000000000000",8408 => "0000000000000000",
8409 => "0000000000000000",8410 => "0000000000000000",
8411 => "0000000000000000",8412 => "0000000000000000",
8413 => "0000000000000000",8414 => "0000000000000000",
8415 => "0000000000000000",8416 => "0000000000000000",
8417 => "0000000000000000",8418 => "0000000000000000",
8419 => "0000000000000000",8420 => "0000000000000000",
8421 => "0000000000000000",8422 => "0000000000000000",
8423 => "0000000000000000",8424 => "0000000000000000",
8425 => "0000000000000000",8426 => "0000000000000000",
8427 => "0000000000000000",8428 => "0000000000000000",
8429 => "0000000000000000",8430 => "0000000000000000",
8431 => "0000000000000000",8432 => "0000000000000000",
8433 => "0000000000000000",8434 => "0000000000000000",
8435 => "0000000000000000",8436 => "0000000000000000",
8437 => "0000000000000000",8438 => "0000000000000000",
8439 => "0000000000000000",8440 => "0000000000000000",
8441 => "0000000000000000",8442 => "0000000000000000",
8443 => "0000000000000000",8444 => "0000000000000000",
8445 => "0000000000000000",8446 => "0000000000000000",
8447 => "0000000000000000",8448 => "0000000000000000",
8449 => "0000000000000000",8450 => "0000000000000000",
8451 => "0000000000000000",8452 => "0000000000000000",
8453 => "0000000000000000",8454 => "0000000000000000",
8455 => "0000000000000000",8456 => "0000000000000000",
8457 => "0000000000000000",8458 => "0000000000000000",
8459 => "0000000000000000",8460 => "0000000000000000",
8461 => "0000000000000000",8462 => "0000000000000000",
8463 => "0000000000000000",8464 => "0000000000000000",
8465 => "0000000000000000",8466 => "0000000000000000",
8467 => "0000000000000000",8468 => "0000000000000000",
8469 => "0000000000000000",8470 => "0000000000000000",
8471 => "0000000000000000",8472 => "0000000000000000",
8473 => "0000000000000000",8474 => "0000000000000000",
8475 => "0000000000000000",8476 => "0000000000000000",
8477 => "0000000000000000",8478 => "0000000000000000",
8479 => "0000000000000000",8480 => "0000000000000000",
8481 => "0000000000000000",8482 => "0000000000000000",
8483 => "0000000000000000",8484 => "0000000000000000",
8485 => "0000000000000000",8486 => "0000000000000000",
8487 => "0000000000000000",8488 => "0000000000000000",
8489 => "0000000000000000",8490 => "0000000000000000",
8491 => "0000000000000000",8492 => "0000000000000000",
8493 => "0000000000000000",8494 => "0000000000000000",
8495 => "0000000000000000",8496 => "0000000000000000",
8497 => "0000000000000000",8498 => "0000000000000000",
8499 => "0000000000000000",8500 => "0000000000000000",
8501 => "0000000000000000",8502 => "0000000000000000",
8503 => "0000000000000000",8504 => "0000000000000000",
8505 => "0000000000000000",8506 => "0000000000000000",
8507 => "0000000000000000",8508 => "0000000000000000",
8509 => "0000000000000000",8510 => "0000000000000000",
8511 => "0000000000000000",8512 => "0000000000000000",
8513 => "0000000000000000",8514 => "0000000000000000",
8515 => "0000000000000000",8516 => "0000000000000000",
8517 => "0000000000000000",8518 => "0000000000000000",
8519 => "0000000000000000",8520 => "0000000000000000",
8521 => "0000000000000000",8522 => "0000000000000000",
8523 => "0000000000000000",8524 => "0000000000000000",
8525 => "0000000000000000",8526 => "0000000000000000",
8527 => "0000000000000000",8528 => "0000000000000000",
8529 => "0000000000000000",8530 => "0000000000000000",
8531 => "0000000000000000",8532 => "0000000000000000",
8533 => "0000000000000000",8534 => "0000000000000000",
8535 => "0000000000000000",8536 => "0000000000000000",
8537 => "0000000000000000",8538 => "0000000000000000",
8539 => "0000000000000000",8540 => "0000000000000000",
8541 => "0000000000000000",8542 => "0000000000000000",
8543 => "0000000000000000",8544 => "0000000000000000",
8545 => "0000000000000000",8546 => "0000000000000000",
8547 => "0000000000000000",8548 => "0000000000000000",
8549 => "0000000000000000",8550 => "0000000000000000",
8551 => "0000000000000000",8552 => "0000000000000000",
8553 => "0000000000000000",8554 => "0000000000000000",
8555 => "0000000000000000",8556 => "0000000000000000",
8557 => "0000000000000000",8558 => "0000000000000000",
8559 => "0000000000000000",8560 => "0000000000000000",
8561 => "0000000000000000",8562 => "0000000000000000",
8563 => "0000000000000000",8564 => "0000000000000000",
8565 => "0000000000000000",8566 => "0000000000000000",
8567 => "0000000000000000",8568 => "0000000000000000",
8569 => "0000000000000000",8570 => "0000000000000000",
8571 => "0000000000000000",8572 => "0000000000000000",
8573 => "0000000000000000",8574 => "0000000000000000",
8575 => "0000000000000000",8576 => "0000000000000000",
8577 => "0000000000000000",8578 => "0000000000000000",
8579 => "0000000000000000",8580 => "0000000000000000",
8581 => "0000000000000000",8582 => "0000000000000000",
8583 => "0000000000000000",8584 => "0000000000000000",
8585 => "0000000000000000",8586 => "0000000000000000",
8587 => "0000000000000000",8588 => "0000000000000000",
8589 => "0000000000000000",8590 => "0000000000000000",
8591 => "0000000000000000",8592 => "0000000000000000",
8593 => "0000000000000000",8594 => "0000000000000000",
8595 => "0000000000000000",8596 => "0000000000000000",
8597 => "0000000000000000",8598 => "0000000000000000",
8599 => "0000000000000000",8600 => "0000000000000000",
8601 => "0000000000000000",8602 => "0000000000000000",
8603 => "0000000000000000",8604 => "0000000000000000",
8605 => "0000000000000000",8606 => "0000000000000000",
8607 => "0000000000000000",8608 => "0000000000000000",
8609 => "0000000000000000",8610 => "0000000000000000",
8611 => "0000000000000000",8612 => "0000000000000000",
8613 => "0000000000000000",8614 => "0000000000000000",
8615 => "0000000000000000",8616 => "0000000000000000",
8617 => "0000000000000000",8618 => "0000000000000000",
8619 => "0000000000000000",8620 => "0000000000000000",
8621 => "0000000000000000",8622 => "0000000000000000",
8623 => "0000000000000000",8624 => "0000000000000000",
8625 => "0000000000000000",8626 => "0000000000000000",
8627 => "0000000000000000",8628 => "0000000000000000",
8629 => "0000000000000000",8630 => "0000000000000000",
8631 => "0000000000000000",8632 => "0000000000000000",
8633 => "0000000000000000",8634 => "0000000000000000",
8635 => "0000000000000000",8636 => "0000000000000000",
8637 => "0000000000000000",8638 => "0000000000000000",
8639 => "0000000000000000",8640 => "0000000000000000",
8641 => "0000000000000000",8642 => "0000000000000000",
8643 => "0000000000000000",8644 => "0000000000000000",
8645 => "0000000000000000",8646 => "0000000000000000",
8647 => "0000000000000000",8648 => "0000000000000000",
8649 => "0000000000000000",8650 => "0000000000000000",
8651 => "0000000000000000",8652 => "0000000000000000",
8653 => "0000000000000000",8654 => "0000000000000000",
8655 => "0000000000000000",8656 => "0000000000000000",
8657 => "0000000000000000",8658 => "0000000000000000",
8659 => "0000000000000000",8660 => "0000000000000000",
8661 => "0000000000000000",8662 => "0000000000000000",
8663 => "0000000000000000",8664 => "0000000000000000",
8665 => "0000000000000000",8666 => "0000000000000000",
8667 => "0000000000000000",8668 => "0000000000000000",
8669 => "0000000000000000",8670 => "0000000000000000",
8671 => "0000000000000000",8672 => "0000000000000000",
8673 => "0000000000000000",8674 => "0000000000000000",
8675 => "0000000000000000",8676 => "0000000000000000",
8677 => "0000000000000000",8678 => "0000000000000000",
8679 => "0000000000000000",8680 => "0000000000000000",
8681 => "0000000000000000",8682 => "0000000000000000",
8683 => "0000000000000000",8684 => "0000000000000000",
8685 => "0000000000000000",8686 => "0000000000000000",
8687 => "0000000000000000",8688 => "0000000000000000",
8689 => "0000000000000000",8690 => "0000000000000000",
8691 => "0000000000000000",8692 => "0000000000000000",
8693 => "0000000000000000",8694 => "0000000000000000",
8695 => "0000000000000000",8696 => "0000000000000000",
8697 => "0000000000000000",8698 => "0000000000000000",
8699 => "0000000000000000",8700 => "0000000000000000",
8701 => "0000000000000000",8702 => "0000000000000000",
8703 => "0000000000000000",8704 => "0000000000000000",
8705 => "0000000000000000",8706 => "0000000000000000",
8707 => "0000000000000000",8708 => "0000000000000000",
8709 => "0000000000000000",8710 => "0000000000000000",
8711 => "0000000000000000",8712 => "0000000000000000",
8713 => "0000000000000000",8714 => "0000000000000000",
8715 => "0000000000000000",8716 => "0000000000000000",
8717 => "0000000000000000",8718 => "0000000000000000",
8719 => "0000000000000000",8720 => "0000000000000000",
8721 => "0000000000000000",8722 => "0000000000000000",
8723 => "0000000000000000",8724 => "0000000000000000",
8725 => "0000000000000000",8726 => "0000000000000000",
8727 => "0000000000000000",8728 => "0000000000000000",
8729 => "0000000000000000",8730 => "0000000000000000",
8731 => "0000000000000000",8732 => "0000000000000000",
8733 => "0000000000000000",8734 => "0000000000000000",
8735 => "0000000000000000",8736 => "0000000000000000",
8737 => "0000000000000000",8738 => "0000000000000000",
8739 => "0000000000000000",8740 => "0000000000000000",
8741 => "0000000000000000",8742 => "0000000000000000",
8743 => "0000000000000000",8744 => "0000000000000000",
8745 => "0000000000000000",8746 => "0000000000000000",
8747 => "0000000000000000",8748 => "0000000000000000",
8749 => "0000000000000000",8750 => "0000000000000000",
8751 => "0000000000000000",8752 => "0000000000000000",
8753 => "0000000000000000",8754 => "0000000000000000",
8755 => "0000000000000000",8756 => "0000000000000000",
8757 => "0000000000000000",8758 => "0000000000000000",
8759 => "0000000000000000",8760 => "0000000000000000",
8761 => "0000000000000000",8762 => "0000000000000000",
8763 => "0000000000000000",8764 => "0000000000000000",
8765 => "0000000000000000",8766 => "0000000000000000",
8767 => "0000000000000000",8768 => "0000000000000000",
8769 => "0000000000000000",8770 => "0000000000000000",
8771 => "0000000000000000",8772 => "0000000000000000",
8773 => "0000000000000000",8774 => "0000000000000000",
8775 => "0000000000000000",8776 => "0000000000000000",
8777 => "0000000000000000",8778 => "0000000000000000",
8779 => "0000000000000000",8780 => "0000000000000000",
8781 => "0000000000000000",8782 => "0000000000000000",
8783 => "0000000000000000",8784 => "0000000000000000",
8785 => "0000000000000000",8786 => "0000000000000000",
8787 => "0000000000000000",8788 => "0000000000000000",
8789 => "0000000000000000",8790 => "0000000000000000",
8791 => "0000000000000000",8792 => "0000000000000000",
8793 => "0000000000000000",8794 => "0000000000000000",
8795 => "0000000000000000",8796 => "0000000000000000",
8797 => "0000000000000000",8798 => "0000000000000000",
8799 => "0000000000000000",8800 => "0000000000000000",
8801 => "0000000000000000",8802 => "0000000000000000",
8803 => "0000000000000000",8804 => "0000000000000000",
8805 => "0000000000000000",8806 => "0000000000000000",
8807 => "0000000000000000",8808 => "0000000000000000",
8809 => "0000000000000000",8810 => "0000000000000000",
8811 => "0000000000000000",8812 => "0000000000000000",
8813 => "0000000000000000",8814 => "0000000000000000",
8815 => "0000000000000000",8816 => "0000000000000000",
8817 => "0000000000000000",8818 => "0000000000000000",
8819 => "0000000000000000",8820 => "0000000000000000",
8821 => "0000000000000000",8822 => "0000000000000000",
8823 => "0000000000000000",8824 => "0000000000000000",
8825 => "0000000000000000",8826 => "0000000000000000",
8827 => "0000000000000000",8828 => "0000000000000000",
8829 => "0000000000000000",8830 => "0000000000000000",
8831 => "0000000000000000",8832 => "0000000000000000",
8833 => "0000000000000000",8834 => "0000000000000000",
8835 => "0000000000000000",8836 => "0000000000000000",
8837 => "0000000000000000",8838 => "0000000000000000",
8839 => "0000000000000000",8840 => "0000000000000000",
8841 => "0000000000000000",8842 => "0000000000000000",
8843 => "0000000000000000",8844 => "0000000000000000",
8845 => "0000000000000000",8846 => "0000000000000000",
8847 => "0000000000000000",8848 => "0000000000000000",
8849 => "0000000000000000",8850 => "0000000000000000",
8851 => "0000000000000000",8852 => "0000000000000000",
8853 => "0000000000000000",8854 => "0000000000000000",
8855 => "0000000000000000",8856 => "0000000000000000",
8857 => "0000000000000000",8858 => "0000000000000000",
8859 => "0000000000000000",8860 => "0000000000000000",
8861 => "0000000000000000",8862 => "0000000000000000",
8863 => "0000000000000000",8864 => "0000000000000000",
8865 => "0000000000000000",8866 => "0000000000000000",
8867 => "0000000000000000",8868 => "0000000000000000",
8869 => "0000000000000000",8870 => "0000000000000000",
8871 => "0000000000000000",8872 => "0000000000000000",
8873 => "0000000000000000",8874 => "0000000000000000",
8875 => "0000000000000000",8876 => "0000000000000000",
8877 => "0000000000000000",8878 => "0000000000000000",
8879 => "0000000000000000",8880 => "0000000000000000",
8881 => "0000000000000000",8882 => "0000000000000000",
8883 => "0000000000000000",8884 => "0000000000000000",
8885 => "0000000000000000",8886 => "0000000000000000",
8887 => "0000000000000000",8888 => "0000000000000000",
8889 => "0000000000000000",8890 => "0000000000000000",
8891 => "0000000000000000",8892 => "0000000000000000",
8893 => "0000000000000000",8894 => "0000000000000000",
8895 => "0000000000000000",8896 => "0000000000000000",
8897 => "0000000000000000",8898 => "0000000000000000",
8899 => "0000000000000000",8900 => "0000000000000000",
8901 => "0000000000000000",8902 => "0000000000000000",
8903 => "0000000000000000",8904 => "0000000000000000",
8905 => "0000000000000000",8906 => "0000000000000000",
8907 => "0000000000000000",8908 => "0000000000000000",
8909 => "0000000000000000",8910 => "0000000000000000",
8911 => "0000000000000000",8912 => "0000000000000000",
8913 => "0000000000000000",8914 => "0000000000000000",
8915 => "0000000000000000",8916 => "0000000000000000",
8917 => "0000000000000000",8918 => "0000000000000000",
8919 => "0000000000000000",8920 => "0000000000000000",
8921 => "0000000000000000",8922 => "0000000000000000",
8923 => "0000000000000000",8924 => "0000000000000000",
8925 => "0000000000000000",8926 => "0000000000000000",
8927 => "0000000000000000",8928 => "0000000000000000",
8929 => "0000000000000000",8930 => "0000000000000000",
8931 => "0000000000000000",8932 => "0000000000000000",
8933 => "0000000000000000",8934 => "0000000000000000",
8935 => "0000000000000000",8936 => "0000000000000000",
8937 => "0000000000000000",8938 => "0000000000000000",
8939 => "0000000000000000",8940 => "0000000000000000",
8941 => "0000000000000000",8942 => "0000000000000000",
8943 => "0000000000000000",8944 => "0000000000000000",
8945 => "0000000000000000",8946 => "0000000000000000",
8947 => "0000000000000000",8948 => "0000000000000000",
8949 => "0000000000000000",8950 => "0000000000000000",
8951 => "0000000000000000",8952 => "0000000000000000",
8953 => "0000000000000000",8954 => "0000000000000000",
8955 => "0000000000000000",8956 => "0000000000000000",
8957 => "0000000000000000",8958 => "0000000000000000",
8959 => "0000000000000000",8960 => "0000000000000000",
8961 => "0000000000000000",8962 => "0000000000000000",
8963 => "0000000000000000",8964 => "0000000000000000",
8965 => "0000000000000000",8966 => "0000000000000000",
8967 => "0000000000000000",8968 => "0000000000000000",
8969 => "0000000000000000",8970 => "0000000000000000",
8971 => "0000000000000000",8972 => "0000000000000000",
8973 => "0000000000000000",8974 => "0000000000000000",
8975 => "0000000000000000",8976 => "0000000000000000",
8977 => "0000000000000000",8978 => "0000000000000000",
8979 => "0000000000000000",8980 => "0000000000000000",
8981 => "0000000000000000",8982 => "0000000000000000",
8983 => "0000000000000000",8984 => "0000000000000000",
8985 => "0000000000000000",8986 => "0000000000000000",
8987 => "0000000000000000",8988 => "0000000000000000",
8989 => "0000000000000000",8990 => "0000000000000000",
8991 => "0000000000000000",8992 => "0000000000000000",
8993 => "0000000000000000",8994 => "0000000000000000",
8995 => "0000000000000000",8996 => "0000000000000000",
8997 => "0000000000000000",8998 => "0000000000000000",
8999 => "0000000000000000",9000 => "0000000000000000",
9001 => "0000000000000000",9002 => "0000000000000000",
9003 => "0000000000000000",9004 => "0000000000000000",
9005 => "0000000000000000",9006 => "0000000000000000",
9007 => "0000000000000000",9008 => "0000000000000000",
9009 => "0000000000000000",9010 => "0000000000000000",
9011 => "0000000000000000",9012 => "0000000000000000",
9013 => "0000000000000000",9014 => "0000000000000000",
9015 => "0000000000000000",9016 => "0000000000000000",
9017 => "0000000000000000",9018 => "0000000000000000",
9019 => "0000000000000000",9020 => "0000000000000000",
9021 => "0000000000000000",9022 => "0000000000000000",
9023 => "0000000000000000",9024 => "0000000000000000",
9025 => "0000000000000000",9026 => "0000000000000000",
9027 => "0000000000000000",9028 => "0000000000000000",
9029 => "0000000000000000",9030 => "0000000000000000",
9031 => "0000000000000000",9032 => "0000000000000000",
9033 => "0000000000000000",9034 => "0000000000000000",
9035 => "0000000000000000",9036 => "0000000000000000",
9037 => "0000000000000000",9038 => "0000000000000000",
9039 => "0000000000000000",9040 => "0000000000000000",
9041 => "0000000000000000",9042 => "0000000000000000",
9043 => "0000000000000000",9044 => "0000000000000000",
9045 => "0000000000000000",9046 => "0000000000000000",
9047 => "0000000000000000",9048 => "0000000000000000",
9049 => "0000000000000000",9050 => "0000000000000000",
9051 => "0000000000000000",9052 => "0000000000000000",
9053 => "0000000000000000",9054 => "0000000000000000",
9055 => "0000000000000000",9056 => "0000000000000000",
9057 => "0000000000000000",9058 => "0000000000000000",
9059 => "0000000000000000",9060 => "0000000000000000",
9061 => "0000000000000000",9062 => "0000000000000000",
9063 => "0000000000000000",9064 => "0000000000000000",
9065 => "0000000000000000",9066 => "0000000000000000",
9067 => "0000000000000000",9068 => "0000000000000000",
9069 => "0000000000000000",9070 => "0000000000000000",
9071 => "0000000000000000",9072 => "0000000000000000",
9073 => "0000000000000000",9074 => "0000000000000000",
9075 => "0000000000000000",9076 => "0000000000000000",
9077 => "0000000000000000",9078 => "0000000000000000",
9079 => "0000000000000000",9080 => "0000000000000000",
9081 => "0000000000000000",9082 => "0000000000000000",
9083 => "0000000000000000",9084 => "0000000000000000",
9085 => "0000000000000000",9086 => "0000000000000000",
9087 => "0000000000000000",9088 => "0000000000000000",
9089 => "0000000000000000",9090 => "0000000000000000",
9091 => "0000000000000000",9092 => "0000000000000000",
9093 => "0000000000000000",9094 => "0000000000000000",
9095 => "0000000000000000",9096 => "0000000000000000",
9097 => "0000000000000000",9098 => "0000000000000000",
9099 => "0000000000000000",9100 => "0000000000000000",
9101 => "0000000000000000",9102 => "0000000000000000",
9103 => "0000000000000000",9104 => "0000000000000000",
9105 => "0000000000000000",9106 => "0000000000000000",
9107 => "0000000000000000",9108 => "0000000000000000",
9109 => "0000000000000000",9110 => "0000000000000000",
9111 => "0000000000000000",9112 => "0000000000000000",
9113 => "0000000000000000",9114 => "0000000000000000",
9115 => "0000000000000000",9116 => "0000000000000000",
9117 => "0000000000000000",9118 => "0000000000000000",
9119 => "0000000000000000",9120 => "0000000000000000",
9121 => "0000000000000000",9122 => "0000000000000000",
9123 => "0000000000000000",9124 => "0000000000000000",
9125 => "0000000000000000",9126 => "0000000000000000",
9127 => "0000000000000000",9128 => "0000000000000000",
9129 => "0000000000000000",9130 => "0000000000000000",
9131 => "0000000000000000",9132 => "0000000000000000",
9133 => "0000000000000000",9134 => "0000000000000000",
9135 => "0000000000000000",9136 => "0000000000000000",
9137 => "0000000000000000",9138 => "0000000000000000",
9139 => "0000000000000000",9140 => "0000000000000000",
9141 => "0000000000000000",9142 => "0000000000000000",
9143 => "0000000000000000",9144 => "0000000000000000",
9145 => "0000000000000000",9146 => "0000000000000000",
9147 => "0000000000000000",9148 => "0000000000000000",
9149 => "0000000000000000",9150 => "0000000000000000",
9151 => "0000000000000000",9152 => "0000000000000000",
9153 => "0000000000000000",9154 => "0000000000000000",
9155 => "0000000000000000",9156 => "0000000000000000",
9157 => "0000000000000000",9158 => "0000000000000000",
9159 => "0000000000000000",9160 => "0000000000000000",
9161 => "0000000000000000",9162 => "0000000000000000",
9163 => "0000000000000000",9164 => "0000000000000000",
9165 => "0000000000000000",9166 => "0000000000000000",
9167 => "0000000000000000",9168 => "0000000000000000",
9169 => "0000000000000000",9170 => "0000000000000000",
9171 => "0000000000000000",9172 => "0000000000000000",
9173 => "0000000000000000",9174 => "0000000000000000",
9175 => "0000000000000000",9176 => "0000000000000000",
9177 => "0000000000000000",9178 => "0000000000000000",
9179 => "0000000000000000",9180 => "0000000000000000",
9181 => "0000000000000000",9182 => "0000000000000000",
9183 => "0000000000000000",9184 => "0000000000000000",
9185 => "0000000000000000",9186 => "0000000000000000",
9187 => "0000000000000000",9188 => "0000000000000000",
9189 => "0000000000000000",9190 => "0000000000000000",
9191 => "0000000000000000",9192 => "0000000000000000",
9193 => "0000000000000000",9194 => "0000000000000000",
9195 => "0000000000000000",9196 => "0000000000000000",
9197 => "0000000000000000",9198 => "0000000000000000",
9199 => "0000000000000000",9200 => "0000000000000000",
9201 => "0000000000000000",9202 => "0000000000000000",
9203 => "0000000000000000",9204 => "0000000000000000",
9205 => "0000000000000000",9206 => "0000000000000000",
9207 => "0000000000000000",9208 => "0000000000000000",
9209 => "0000000000000000",9210 => "0000000000000000",
9211 => "0000000000000000",9212 => "0000000000000000",
9213 => "0000000000000000",9214 => "0000000000000000",
9215 => "0000000000000000",9216 => "0000000000000000",
9217 => "0000000000000000",9218 => "0000000000000000",
9219 => "0000000000000000",9220 => "0000000000000000",
9221 => "0000000000000000",9222 => "0000000000000000",
9223 => "0000000000000000",9224 => "0000000000000000",
9225 => "0000000000000000",9226 => "0000000000000000",
9227 => "0000000000000000",9228 => "0000000000000000",
9229 => "0000000000000000",9230 => "0000000000000000",
9231 => "0000000000000000",9232 => "0000000000000000",
9233 => "0000000000000000",9234 => "0000000000000000",
9235 => "0000000000000000",9236 => "0000000000000000",
9237 => "0000000000000000",9238 => "0000000000000000",
9239 => "0000000000000000",9240 => "0000000000000000",
9241 => "0000000000000000",9242 => "0000000000000000",
9243 => "0000000000000000",9244 => "0000000000000000",
9245 => "0000000000000000",9246 => "0000000000000000",
9247 => "0000000000000000",9248 => "0000000000000000",
9249 => "0000000000000000",9250 => "0000000000000000",
9251 => "0000000000000000",9252 => "0000000000000000",
9253 => "0000000000000000",9254 => "0000000000000000",
9255 => "0000000000000000",9256 => "0000000000000000",
9257 => "0000000000000000",9258 => "0000000000000000",
9259 => "0000000000000000",9260 => "0000000000000000",
9261 => "0000000000000000",9262 => "0000000000000000",
9263 => "0000000000000000",9264 => "0000000000000000",
9265 => "0000000000000000",9266 => "0000000000000000",
9267 => "0000000000000000",9268 => "0000000000000000",
9269 => "0000000000000000",9270 => "0000000000000000",
9271 => "0000000000000000",9272 => "0000000000000000",
9273 => "0000000000000000",9274 => "0000000000000000",
9275 => "0000000000000000",9276 => "0000000000000000",
9277 => "0000000000000000",9278 => "0000000000000000",
9279 => "0000000000000000",9280 => "0000000000000000",
9281 => "0000000000000000",9282 => "0000000000000000",
9283 => "0000000000000000",9284 => "0000000000000000",
9285 => "0000000000000000",9286 => "0000000000000000",
9287 => "0000000000000000",9288 => "0000000000000000",
9289 => "0000000000000000",9290 => "0000000000000000",
9291 => "0000000000000000",9292 => "0000000000000000",
9293 => "0000000000000000",9294 => "0000000000000000",
9295 => "0000000000000000",9296 => "0000000000000000",
9297 => "0000000000000000",9298 => "0000000000000000",
9299 => "0000000000000000",9300 => "0000000000000000",
9301 => "0000000000000000",9302 => "0000000000000000",
9303 => "0000000000000000",9304 => "0000000000000000",
9305 => "0000000000000000",9306 => "0000000000000000",
9307 => "0000000000000000",9308 => "0000000000000000",
9309 => "0000000000000000",9310 => "0000000000000000",
9311 => "0000000000000000",9312 => "0000000000000000",
9313 => "0000000000000000",9314 => "0000000000000000",
9315 => "0000000000000000",9316 => "0000000000000000",
9317 => "0000000000000000",9318 => "0000000000000000",
9319 => "0000000000000000",9320 => "0000000000000000",
9321 => "0000000000000000",9322 => "0000000000000000",
9323 => "0000000000000000",9324 => "0000000000000000",
9325 => "0000000000000000",9326 => "0000000000000000",
9327 => "0000000000000000",9328 => "0000000000000000",
9329 => "0000000000000000",9330 => "0000000000000000",
9331 => "0000000000000000",9332 => "0000000000000000",
9333 => "0000000000000000",9334 => "0000000000000000",
9335 => "0000000000000000",9336 => "0000000000000000",
9337 => "0000000000000000",9338 => "0000000000000000",
9339 => "0000000000000000",9340 => "0000000000000000",
9341 => "0000000000000000",9342 => "0000000000000000",
9343 => "0000000000000000",9344 => "0000000000000000",
9345 => "0000000000000000",9346 => "0000000000000000",
9347 => "0000000000000000",9348 => "0000000000000000",
9349 => "0000000000000000",9350 => "0000000000000000",
9351 => "0000000000000000",9352 => "0000000000000000",
9353 => "0000000000000000",9354 => "0000000000000000",
9355 => "0000000000000000",9356 => "0000000000000000",
9357 => "0000000000000000",9358 => "0000000000000000",
9359 => "0000000000000000",9360 => "0000000000000000",
9361 => "0000000000000000",9362 => "0000000000000000",
9363 => "0000000000000000",9364 => "0000000000000000",
9365 => "0000000000000000",9366 => "0000000000000000",
9367 => "0000000000000000",9368 => "0000000000000000",
9369 => "0000000000000000",9370 => "0000000000000000",
9371 => "0000000000000000",9372 => "0000000000000000",
9373 => "0000000000000000",9374 => "0000000000000000",
9375 => "0000000000000000",9376 => "0000000000000000",
9377 => "0000000000000000",9378 => "0000000000000000",
9379 => "0000000000000000",9380 => "0000000000000000",
9381 => "0000000000000000",9382 => "0000000000000000",
9383 => "0000000000000000",9384 => "0000000000000000",
9385 => "0000000000000000",9386 => "0000000000000000",
9387 => "0000000000000000",9388 => "0000000000000000",
9389 => "0000000000000000",9390 => "0000000000000000",
9391 => "0000000000000000",9392 => "0000000000000000",
9393 => "0000000000000000",9394 => "0000000000000000",
9395 => "0000000000000000",9396 => "0000000000000000",
9397 => "0000000000000000",9398 => "0000000000000000",
9399 => "0000000000000000",9400 => "0000000000000000",
9401 => "0000000000000000",9402 => "0000000000000000",
9403 => "0000000000000000",9404 => "0000000000000000",
9405 => "0000000000000000",9406 => "0000000000000000",
9407 => "0000000000000000",9408 => "0000000000000000",
9409 => "0000000000000000",9410 => "0000000000000000",
9411 => "0000000000000000",9412 => "0000000000000000",
9413 => "0000000000000000",9414 => "0000000000000000",
9415 => "0000000000000000",9416 => "0000000000000000",
9417 => "0000000000000000",9418 => "0000000000000000",
9419 => "0000000000000000",9420 => "0000000000000000",
9421 => "0000000000000000",9422 => "0000000000000000",
9423 => "0000000000000000",9424 => "0000000000000000",
9425 => "0000000000000000",9426 => "0000000000000000",
9427 => "0000000000000000",9428 => "0000000000000000",
9429 => "0000000000000000",9430 => "0000000000000000",
9431 => "0000000000000000",9432 => "0000000000000000",
9433 => "0000000000000000",9434 => "0000000000000000",
9435 => "0000000000000000",9436 => "0000000000000000",
9437 => "0000000000000000",9438 => "0000000000000000",
9439 => "0000000000000000",9440 => "0000000000000000",
9441 => "0000000000000000",9442 => "0000000000000000",
9443 => "0000000000000000",9444 => "0000000000000000",
9445 => "0000000000000000",9446 => "0000000000000000",
9447 => "0000000000000000",9448 => "0000000000000000",
9449 => "0000000000000000",9450 => "0000000000000000",
9451 => "0000000000000000",9452 => "0000000000000000",
9453 => "0000000000000000",9454 => "0000000000000000",
9455 => "0000000000000000",9456 => "0000000000000000",
9457 => "0000000000000000",9458 => "0000000000000000",
9459 => "0000000000000000",9460 => "0000000000000000",
9461 => "0000000000000000",9462 => "0000000000000000",
9463 => "0000000000000000",9464 => "0000000000000000",
9465 => "0000000000000000",9466 => "0000000000000000",
9467 => "0000000000000000",9468 => "0000000000000000",
9469 => "0000000000000000",9470 => "0000000000000000",
9471 => "0000000000000000",9472 => "0000000000000000",
9473 => "0000000000000000",9474 => "0000000000000000",
9475 => "0000000000000000",9476 => "0000000000000000",
9477 => "0000000000000000",9478 => "0000000000000000",
9479 => "0000000000000000",9480 => "0000000000000000",
9481 => "0000000000000000",9482 => "0000000000000000",
9483 => "0000000000000000",9484 => "0000000000000000",
9485 => "0000000000000000",9486 => "0000000000000000",
9487 => "0000000000000000",9488 => "0000000000000000",
9489 => "0000000000000000",9490 => "0000000000000000",
9491 => "0000000000000000",9492 => "0000000000000000",
9493 => "0000000000000000",9494 => "0000000000000000",
9495 => "0000000000000000",9496 => "0000000000000000",
9497 => "0000000000000000",9498 => "0000000000000000",
9499 => "0000000000000000",9500 => "0000000000000000",
9501 => "0000000000000000",9502 => "0000000000000000",
9503 => "0000000000000000",9504 => "0000000000000000",
9505 => "0000000000000000",9506 => "0000000000000000",
9507 => "0000000000000000",9508 => "0000000000000000",
9509 => "0000000000000000",9510 => "0000000000000000",
9511 => "0000000000000000",9512 => "0000000000000000",
9513 => "0000000000000000",9514 => "0000000000000000",
9515 => "0000000000000000",9516 => "0000000000000000",
9517 => "0000000000000000",9518 => "0000000000000000",
9519 => "0000000000000000",9520 => "0000000000000000",
9521 => "0000000000000000",9522 => "0000000000000000",
9523 => "0000000000000000",9524 => "0000000000000000",
9525 => "0000000000000000",9526 => "0000000000000000",
9527 => "0000000000000000",9528 => "0000000000000000",
9529 => "0000000000000000",9530 => "0000000000000000",
9531 => "0000000000000000",9532 => "0000000000000000",
9533 => "0000000000000000",9534 => "0000000000000000",
9535 => "0000000000000000",9536 => "0000000000000000",
9537 => "0000000000000000",9538 => "0000000000000000",
9539 => "0000000000000000",9540 => "0000000000000000",
9541 => "0000000000000000",9542 => "0000000000000000",
9543 => "0000000000000000",9544 => "0000000000000000",
9545 => "0000000000000000",9546 => "0000000000000000",
9547 => "0000000000000000",9548 => "0000000000000000",
9549 => "0000000000000000",9550 => "0000000000000000",
9551 => "0000000000000000",9552 => "0000000000000000",
9553 => "0000000000000000",9554 => "0000000000000000",
9555 => "0000000000000000",9556 => "0000000000000000",
9557 => "0000000000000000",9558 => "0000000000000000",
9559 => "0000000000000000",9560 => "0000000000000000",
9561 => "0000000000000000",9562 => "0000000000000000",
9563 => "0000000000000000",9564 => "0000000000000000",
9565 => "0000000000000000",9566 => "0000000000000000",
9567 => "0000000000000000",9568 => "0000000000000000",
9569 => "0000000000000000",9570 => "0000000000000000",
9571 => "0000000000000000",9572 => "0000000000000000",
9573 => "0000000000000000",9574 => "0000000000000000",
9575 => "0000000000000000",9576 => "0000000000000000",
9577 => "0000000000000000",9578 => "0000000000000000",
9579 => "0000000000000000",9580 => "0000000000000000",
9581 => "0000000000000000",9582 => "0000000000000000",
9583 => "0000000000000000",9584 => "0000000000000000",
9585 => "0000000000000000",9586 => "0000000000000000",
9587 => "0000000000000000",9588 => "0000000000000000",
9589 => "0000000000000000",9590 => "0000000000000000",
9591 => "0000000000000000",9592 => "0000000000000000",
9593 => "0000000000000000",9594 => "0000000000000000",
9595 => "0000000000000000",9596 => "0000000000000000",
9597 => "0000000000000000",9598 => "0000000000000000",
9599 => "0000000000000000",9600 => "0000000000000000",
9601 => "0000000000000000",9602 => "0000000000000000",
9603 => "0000000000000000",9604 => "0000000000000000",
9605 => "0000000000000000",9606 => "0000000000000000",
9607 => "0000000000000000",9608 => "0000000000000000",
9609 => "0000000000000000",9610 => "0000000000000000",
9611 => "0000000000000000",9612 => "0000000000000000",
9613 => "0000000000000000",9614 => "0000000000000000",
9615 => "0000000000000000",9616 => "0000000000000000",
9617 => "0000000000000000",9618 => "0000000000000000",
9619 => "0000000000000000",9620 => "0000000000000000",
9621 => "0000000000000000",9622 => "0000000000000000",
9623 => "0000000000000000",9624 => "0000000000000000",
9625 => "0000000000000000",9626 => "0000000000000000",
9627 => "0000000000000000",9628 => "0000000000000000",
9629 => "0000000000000000",9630 => "0000000000000000",
9631 => "0000000000000000",9632 => "0000000000000000",
9633 => "0000000000000000",9634 => "0000000000000000",
9635 => "0000000000000000",9636 => "0000000000000000",
9637 => "0000000000000000",9638 => "0000000000000000",
9639 => "0000000000000000",9640 => "0000000000000000",
9641 => "0000000000000000",9642 => "0000000000000000",
9643 => "0000000000000000",9644 => "0000000000000000",
9645 => "0000000000000000",9646 => "0000000000000000",
9647 => "0000000000000000",9648 => "0000000000000000",
9649 => "0000000000000000",9650 => "0000000000000000",
9651 => "0000000000000000",9652 => "0000000000000000",
9653 => "0000000000000000",9654 => "0000000000000000",
9655 => "0000000000000000",9656 => "0000000000000000",
9657 => "0000000000000000",9658 => "0000000000000000",
9659 => "0000000000000000",9660 => "0000000000000000",
9661 => "0000000000000000",9662 => "0000000000000000",
9663 => "0000000000000000",9664 => "0000000000000000",
9665 => "0000000000000000",9666 => "0000000000000000",
9667 => "0000000000000000",9668 => "0000000000000000",
9669 => "0000000000000000",9670 => "0000000000000000",
9671 => "0000000000000000",9672 => "0000000000000000",
9673 => "0000000000000000",9674 => "0000000000000000",
9675 => "0000000000000000",9676 => "0000000000000000",
9677 => "0000000000000000",9678 => "0000000000000000",
9679 => "0000000000000000",9680 => "0000000000000000",
9681 => "0000000000000000",9682 => "0000000000000000",
9683 => "0000000000000000",9684 => "0000000000000000",
9685 => "0000000000000000",9686 => "0000000000000000",
9687 => "0000000000000000",9688 => "0000000000000000",
9689 => "0000000000000000",9690 => "0000000000000000",
9691 => "0000000000000000",9692 => "0000000000000000",
9693 => "0000000000000000",9694 => "0000000000000000",
9695 => "0000000000000000",9696 => "0000000000000000",
9697 => "0000000000000000",9698 => "0000000000000000",
9699 => "0000000000000000",9700 => "0000000000000000",
9701 => "0000000000000000",9702 => "0000000000000000",
9703 => "0000000000000000",9704 => "0000000000000000",
9705 => "0000000000000000",9706 => "0000000000000000",
9707 => "0000000000000000",9708 => "0000000000000000",
9709 => "0000000000000000",9710 => "0000000000000000",
9711 => "0000000000000000",9712 => "0000000000000000",
9713 => "0000000000000000",9714 => "0000000000000000",
9715 => "0000000000000000",9716 => "0000000000000000",
9717 => "0000000000000000",9718 => "0000000000000000",
9719 => "0000000000000000",9720 => "0000000000000000",
9721 => "0000000000000000",9722 => "0000000000000000",
9723 => "0000000000000000",9724 => "0000000000000000",
9725 => "0000000000000000",9726 => "0000000000000000",
9727 => "0000000000000000",9728 => "0000000000000000",
9729 => "0000000000000000",9730 => "0000000000000000",
9731 => "0000000000000000",9732 => "0000000000000000",
9733 => "0000000000000000",9734 => "0000000000000000",
9735 => "0000000000000000",9736 => "0000000000000000",
9737 => "0000000000000000",9738 => "0000000000000000",
9739 => "0000000000000000",9740 => "0000000000000000",
9741 => "0000000000000000",9742 => "0000000000000000",
9743 => "0000000000000000",9744 => "0000000000000000",
9745 => "0000000000000000",9746 => "0000000000000000",
9747 => "0000000000000000",9748 => "0000000000000000",
9749 => "0000000000000000",9750 => "0000000000000000",
9751 => "0000000000000000",9752 => "0000000000000000",
9753 => "0000000000000000",9754 => "0000000000000000",
9755 => "0000000000000000",9756 => "0000000000000000",
9757 => "0000000000000000",9758 => "0000000000000000",
9759 => "0000000000000000",9760 => "0000000000000000",
9761 => "0000000000000000",9762 => "0000000000000000",
9763 => "0000000000000000",9764 => "0000000000000000",
9765 => "0000000000000000",9766 => "0000000000000000",
9767 => "0000000000000000",9768 => "0000000000000000",
9769 => "0000000000000000",9770 => "0000000000000000",
9771 => "0000000000000000",9772 => "0000000000000000",
9773 => "0000000000000000",9774 => "0000000000000000",
9775 => "0000000000000000",9776 => "0000000000000000",
9777 => "0000000000000000",9778 => "0000000000000000",
9779 => "0000000000000000",9780 => "0000000000000000",
9781 => "0000000000000000",9782 => "0000000000000000",
9783 => "0000000000000000",9784 => "0000000000000000",
9785 => "0000000000000000",9786 => "0000000000000000",
9787 => "0000000000000000",9788 => "0000000000000000",
9789 => "0000000000000000",9790 => "0000000000000000",
9791 => "0000000000000000",9792 => "0000000000000000",
9793 => "0000000000000000",9794 => "0000000000000000",
9795 => "0000000000000000",9796 => "0000000000000000",
9797 => "0000000000000000",9798 => "0000000000000000",
9799 => "0000000000000000",9800 => "0000000000000000",
9801 => "0000000000000000",9802 => "0000000000000000",
9803 => "0000000000000000",9804 => "0000000000000000",
9805 => "0000000000000000",9806 => "0000000000000000",
9807 => "0000000000000000",9808 => "0000000000000000",
9809 => "0000000000000000",9810 => "0000000000000000",
9811 => "0000000000000000",9812 => "0000000000000000",
9813 => "0000000000000000",9814 => "0000000000000000",
9815 => "0000000000000000",9816 => "0000000000000000",
9817 => "0000000000000000",9818 => "0000000000000000",
9819 => "0000000000000000",9820 => "0000000000000000",
9821 => "0000000000000000",9822 => "0000000000000000",
9823 => "0000000000000000",9824 => "0000000000000000",
9825 => "0000000000000000",9826 => "0000000000000000",
9827 => "0000000000000000",9828 => "0000000000000000",
9829 => "0000000000000000",9830 => "0000000000000000",
9831 => "0000000000000000",9832 => "0000000000000000",
9833 => "0000000000000000",9834 => "0000000000000000",
9835 => "0000000000000000",9836 => "0000000000000000",
9837 => "0000000000000000",9838 => "0000000000000000",
9839 => "0000000000000000",9840 => "0000000000000000",
9841 => "0000000000000000",9842 => "0000000000000000",
9843 => "0000000000000000",9844 => "0000000000000000",
9845 => "0000000000000000",9846 => "0000000000000000",
9847 => "0000000000000000",9848 => "0000000000000000",
9849 => "0000000000000000",9850 => "0000000000000000",
9851 => "0000000000000000",9852 => "0000000000000000",
9853 => "0000000000000000",9854 => "0000000000000000",
9855 => "0000000000000000",9856 => "0000000000000000",
9857 => "0000000000000000",9858 => "0000000000000000",
9859 => "0000000000000000",9860 => "0000000000000000",
9861 => "0000000000000000",9862 => "0000000000000000",
9863 => "0000000000000000",9864 => "0000000000000000",
9865 => "0000000000000000",9866 => "0000000000000000",
9867 => "0000000000000000",9868 => "0000000000000000",
9869 => "0000000000000000",9870 => "0000000000000000",
9871 => "0000000000000000",9872 => "0000000000000000",
9873 => "0000000000000000",9874 => "0000000000000000",
9875 => "0000000000000000",9876 => "0000000000000000",
9877 => "0000000000000000",9878 => "0000000000000000",
9879 => "0000000000000000",9880 => "0000000000000000",
9881 => "0000000000000000",9882 => "0000000000000000",
9883 => "0000000000000000",9884 => "0000000000000000",
9885 => "0000000000000000",9886 => "0000000000000000",
9887 => "0000000000000000",9888 => "0000000000000000",
9889 => "0000000000000000",9890 => "0000000000000000",
9891 => "0000000000000000",9892 => "0000000000000000",
9893 => "0000000000000000",9894 => "0000000000000000",
9895 => "0000000000000000",9896 => "0000000000000000",
9897 => "0000000000000000",9898 => "0000000000000000",
9899 => "0000000000000000",9900 => "0000000000000000",
9901 => "0000000000000000",9902 => "0000000000000000",
9903 => "0000000000000000",9904 => "0000000000000000",
9905 => "0000000000000000",9906 => "0000000000000000",
9907 => "0000000000000000",9908 => "0000000000000000",
9909 => "0000000000000000",9910 => "0000000000000000",
9911 => "0000000000000000",9912 => "0000000000000000",
9913 => "0000000000000000",9914 => "0000000000000000",
9915 => "0000000000000000",9916 => "0000000000000000",
9917 => "0000000000000000",9918 => "0000000000000000",
9919 => "0000000000000000",9920 => "0000000000000000",
9921 => "0000000000000000",9922 => "0000000000000000",
9923 => "0000000000000000",9924 => "0000000000000000",
9925 => "0000000000000000",9926 => "0000000000000000",
9927 => "0000000000000000",9928 => "0000000000000000",
9929 => "0000000000000000",9930 => "0000000000000000",
9931 => "0000000000000000",9932 => "0000000000000000",
9933 => "0000000000000000",9934 => "0000000000000000",
9935 => "0000000000000000",9936 => "0000000000000000",
9937 => "0000000000000000",9938 => "0000000000000000",
9939 => "0000000000000000",9940 => "0000000000000000",
9941 => "0000000000000000",9942 => "0000000000000000",
9943 => "0000000000000000",9944 => "0000000000000000",
9945 => "0000000000000000",9946 => "0000000000000000",
9947 => "0000000000000000",9948 => "0000000000000000",
9949 => "0000000000000000",9950 => "0000000000000000",
9951 => "0000000000000000",9952 => "0000000000000000",
9953 => "0000000000000000",9954 => "0000000000000000",
9955 => "0000000000000000",9956 => "0000000000000000",
9957 => "0000000000000000",9958 => "0000000000000000",
9959 => "0000000000000000",9960 => "0000000000000000",
9961 => "0000000000000000",9962 => "0000000000000000",
9963 => "0000000000000000",9964 => "0000000000000000",
9965 => "0000000000000000",9966 => "0000000000000000",
9967 => "0000000000000000",9968 => "0000000000000000",
9969 => "0000000000000000",9970 => "0000000000000000",
9971 => "0000000000000000",9972 => "0000000000000000",
9973 => "0000000000000000",9974 => "0000000000000000",
9975 => "0000000000000000",9976 => "0000000000000000",
9977 => "0000000000000000",9978 => "0000000000000000",
9979 => "0000000000000000",9980 => "0000000000000000",
9981 => "0000000000000000",9982 => "0000000000000000",
9983 => "0000000000000000",9984 => "0000000000000000",
9985 => "0000000000000000",9986 => "0000000000000000",
9987 => "0000000000000000",9988 => "0000000000000000",
9989 => "0000000000000000",9990 => "0000000000000000",
9991 => "0000000000000000",9992 => "0000000000000000",
9993 => "0000000000000000",9994 => "0000000000000000",
9995 => "0000000000000000",9996 => "0000000000000000",
9997 => "0000000000000000",9998 => "0000000000000000",
9999 => "0000000000000000",10000 => "0000000000000000",
10001 => "0000000000000000",10002 => "0000000000000000",
10003 => "0000000000000000",10004 => "0000000000000000",
10005 => "0000000000000000",10006 => "0000000000000000",
10007 => "0000000000000000",10008 => "0000000000000000",
10009 => "0000000000000000",10010 => "0000000000000000",
10011 => "0000000000000000",10012 => "0000000000000000",
10013 => "0000000000000000",10014 => "0000000000000000",
10015 => "0000000000000000",10016 => "0000000000000000",
10017 => "0000000000000000",10018 => "0000000000000000",
10019 => "0000000000000000",10020 => "0000000000000000",
10021 => "0000000000000000",10022 => "0000000000000000",
10023 => "0000000000000000",10024 => "0000000000000000",
10025 => "0000000000000000",10026 => "0000000000000000",
10027 => "0000000000000000",10028 => "0000000000000000",
10029 => "0000000000000000",10030 => "0000000000000000",
10031 => "0000000000000000",10032 => "0000000000000000",
10033 => "0000000000000000",10034 => "0000000000000000",
10035 => "0000000000000000",10036 => "0000000000000000",
10037 => "0000000000000000",10038 => "0000000000000000",
10039 => "0000000000000000",10040 => "0000000000000000",
10041 => "0000000000000000",10042 => "0000000000000000",
10043 => "0000000000000000",10044 => "0000000000000000",
10045 => "0000000000000000",10046 => "0000000000000000",
10047 => "0000000000000000",10048 => "0000000000000000",
10049 => "0000000000000000",10050 => "0000000000000000",
10051 => "0000000000000000",10052 => "0000000000000000",
10053 => "0000000000000000",10054 => "0000000000000000",
10055 => "0000000000000000",10056 => "0000000000000000",
10057 => "0000000000000000",10058 => "0000000000000000",
10059 => "0000000000000000",10060 => "0000000000000000",
10061 => "0000000000000000",10062 => "0000000000000000",
10063 => "0000000000000000",10064 => "0000000000000000",
10065 => "0000000000000000",10066 => "0000000000000000",
10067 => "0000000000000000",10068 => "0000000000000000",
10069 => "0000000000000000",10070 => "0000000000000000",
10071 => "0000000000000000",10072 => "0000000000000000",
10073 => "0000000000000000",10074 => "0000000000000000",
10075 => "0000000000000000",10076 => "0000000000000000",
10077 => "0000000000000000",10078 => "0000000000000000",
10079 => "0000000000000000",10080 => "0000000000000000",
10081 => "0000000000000000",10082 => "0000000000000000",
10083 => "0000000000000000",10084 => "0000000000000000",
10085 => "0000000000000000",10086 => "0000000000000000",
10087 => "0000000000000000",10088 => "0000000000000000",
10089 => "0000000000000000",10090 => "0000000000000000",
10091 => "0000000000000000",10092 => "0000000000000000",
10093 => "0000000000000000",10094 => "0000000000000000",
10095 => "0000000000000000",10096 => "0000000000000000",
10097 => "0000000000000000",10098 => "0000000000000000",
10099 => "0000000000000000",10100 => "0000000000000000",
10101 => "0000000000000000",10102 => "0000000000000000",
10103 => "0000000000000000",10104 => "0000000000000000",
10105 => "0000000000000000",10106 => "0000000000000000",
10107 => "0000000000000000",10108 => "0000000000000000",
10109 => "0000000000000000",10110 => "0000000000000000",
10111 => "0000000000000000",10112 => "0000000000000000",
10113 => "0000000000000000",10114 => "0000000000000000",
10115 => "0000000000000000",10116 => "0000000000000000",
10117 => "0000000000000000",10118 => "0000000000000000",
10119 => "0000000000000000",10120 => "0000000000000000",
10121 => "0000000000000000",10122 => "0000000000000000",
10123 => "0000000000000000",10124 => "0000000000000000",
10125 => "0000000000000000",10126 => "0000000000000000",
10127 => "0000000000000000",10128 => "0000000000000000",
10129 => "0000000000000000",10130 => "0000000000000000",
10131 => "0000000000000000",10132 => "0000000000000000",
10133 => "0000000000000000",10134 => "0000000000000000",
10135 => "0000000000000000",10136 => "0000000000000000",
10137 => "0000000000000000",10138 => "0000000000000000",
10139 => "0000000000000000",10140 => "0000000000000000",
10141 => "0000000000000000",10142 => "0000000000000000",
10143 => "0000000000000000",10144 => "0000000000000000",
10145 => "0000000000000000",10146 => "0000000000000000",
10147 => "0000000000000000",10148 => "0000000000000000",
10149 => "0000000000000000",10150 => "0000000000000000",
10151 => "0000000000000000",10152 => "0000000000000000",
10153 => "0000000000000000",10154 => "0000000000000000",
10155 => "0000000000000000",10156 => "0000000000000000",
10157 => "0000000000000000",10158 => "0000000000000000",
10159 => "0000000000000000",10160 => "0000000000000000",
10161 => "0000000000000000",10162 => "0000000000000000",
10163 => "0000000000000000",10164 => "0000000000000000",
10165 => "0000000000000000",10166 => "0000000000000000",
10167 => "0000000000000000",10168 => "0000000000000000",
10169 => "0000000000000000",10170 => "0000000000000000",
10171 => "0000000000000000",10172 => "0000000000000000",
10173 => "0000000000000000",10174 => "0000000000000000",
10175 => "0000000000000000",10176 => "0000000000000000",
10177 => "0000000000000000",10178 => "0000000000000000",
10179 => "0000000000000000",10180 => "0000000000000000",
10181 => "0000000000000000",10182 => "0000000000000000",
10183 => "0000000000000000",10184 => "0000000000000000",
10185 => "0000000000000000",10186 => "0000000000000000",
10187 => "0000000000000000",10188 => "0000000000000000",
10189 => "0000000000000000",10190 => "0000000000000000",
10191 => "0000000000000000",10192 => "0000000000000000",
10193 => "0000000000000000",10194 => "0000000000000000",
10195 => "0000000000000000",10196 => "0000000000000000",
10197 => "0000000000000000",10198 => "0000000000000000",
10199 => "0000000000000000",10200 => "0000000000000000",
10201 => "0000000000000000",10202 => "0000000000000000",
10203 => "0000000000000000",10204 => "0000000000000000",
10205 => "0000000000000000",10206 => "0000000000000000",
10207 => "0000000000000000",10208 => "0000000000000000",
10209 => "0000000000000000",10210 => "0000000000000000",
10211 => "0000000000000000",10212 => "0000000000000000",
10213 => "0000000000000000",10214 => "0000000000000000",
10215 => "0000000000000000",10216 => "0000000000000000",
10217 => "0000000000000000",10218 => "0000000000000000",
10219 => "0000000000000000",10220 => "0000000000000000",
10221 => "0000000000000000",10222 => "0000000000000000",
10223 => "0000000000000000",10224 => "0000000000000000",
10225 => "0000000000000000",10226 => "0000000000000000",
10227 => "0000000000000000",10228 => "0000000000000000",
10229 => "0000000000000000",10230 => "0000000000000000",
10231 => "0000000000000000",10232 => "0000000000000000",
10233 => "0000000000000000",10234 => "0000000000000000",
10235 => "0000000000000000",10236 => "0000000000000000",
10237 => "0000000000000000",10238 => "0000000000000000",
10239 => "0000000000000000",10240 => "0000000000000000",
10241 => "0000000000000000",10242 => "0000000000000000",
10243 => "0000000000000000",10244 => "0000000000000000",
10245 => "0000000000000000",10246 => "0000000000000000",
10247 => "0000000000000000",10248 => "0000000000000000",
10249 => "0000000000000000",10250 => "0000000000000000",
10251 => "0000000000000000",10252 => "0000000000000000",
10253 => "0000000000000000",10254 => "0000000000000000",
10255 => "0000000000000000",10256 => "0000000000000000",
10257 => "0000000000000000",10258 => "0000000000000000",
10259 => "0000000000000000",10260 => "0000000000000000",
10261 => "0000000000000000",10262 => "0000000000000000",
10263 => "0000000000000000",10264 => "0000000000000000",
10265 => "0000000000000000",10266 => "0000000000000000",
10267 => "0000000000000000",10268 => "0000000000000000",
10269 => "0000000000000000",10270 => "0000000000000000",
10271 => "0000000000000000",10272 => "0000000000000000",
10273 => "0000000000000000",10274 => "0000000000000000",
10275 => "0000000000000000",10276 => "0000000000000000",
10277 => "0000000000000000",10278 => "0000000000000000",
10279 => "0000000000000000",10280 => "0000000000000000",
10281 => "0000000000000000",10282 => "0000000000000000",
10283 => "0000000000000000",10284 => "0000000000000000",
10285 => "0000000000000000",10286 => "0000000000000000",
10287 => "0000000000000000",10288 => "0000000000000000",
10289 => "0000000000000000",10290 => "0000000000000000",
10291 => "0000000000000000",10292 => "0000000000000000",
10293 => "0000000000000000",10294 => "0000000000000000",
10295 => "0000000000000000",10296 => "0000000000000000",
10297 => "0000000000000000",10298 => "0000000000000000",
10299 => "0000000000000000",10300 => "0000000000000000",
10301 => "0000000000000000",10302 => "0000000000000000",
10303 => "0000000000000000",10304 => "0000000000000000",
10305 => "0000000000000000",10306 => "0000000000000000",
10307 => "0000000000000000",10308 => "0000000000000000",
10309 => "0000000000000000",10310 => "0000000000000000",
10311 => "0000000000000000",10312 => "0000000000000000",
10313 => "0000000000000000",10314 => "0000000000000000",
10315 => "0000000000000000",10316 => "0000000000000000",
10317 => "0000000000000000",10318 => "0000000000000000",
10319 => "0000000000000000",10320 => "0000000000000000",
10321 => "0000000000000000",10322 => "0000000000000000",
10323 => "0000000000000000",10324 => "0000000000000000",
10325 => "0000000000000000",10326 => "0000000000000000",
10327 => "0000000000000000",10328 => "0000000000000000",
10329 => "0000000000000000",10330 => "0000000000000000",
10331 => "0000000000000000",10332 => "0000000000000000",
10333 => "0000000000000000",10334 => "0000000000000000",
10335 => "0000000000000000",10336 => "0000000000000000",
10337 => "0000000000000000",10338 => "0000000000000000",
10339 => "0000000000000000",10340 => "0000000000000000",
10341 => "0000000000000000",10342 => "0000000000000000",
10343 => "0000000000000000",10344 => "0000000000000000",
10345 => "0000000000000000",10346 => "0000000000000000",
10347 => "0000000000000000",10348 => "0000000000000000",
10349 => "0000000000000000",10350 => "0000000000000000",
10351 => "0000000000000000",10352 => "0000000000000000",
10353 => "0000000000000000",10354 => "0000000000000000",
10355 => "0000000000000000",10356 => "0000000000000000",
10357 => "0000000000000000",10358 => "0000000000000000",
10359 => "0000000000000000",10360 => "0000000000000000",
10361 => "0000000000000000",10362 => "0000000000000000",
10363 => "0000000000000000",10364 => "0000000000000000",
10365 => "0000000000000000",10366 => "0000000000000000",
10367 => "0000000000000000",10368 => "0000000000000000",
10369 => "0000000000000000",10370 => "0000000000000000",
10371 => "0000000000000000",10372 => "0000000000000000",
10373 => "0000000000000000",10374 => "0000000000000000",
10375 => "0000000000000000",10376 => "0000000000000000",
10377 => "0000000000000000",10378 => "0000000000000000",
10379 => "0000000000000000",10380 => "0000000000000000",
10381 => "0000000000000000",10382 => "0000000000000000",
10383 => "0000000000000000",10384 => "0000000000000000",
10385 => "0000000000000000",10386 => "0000000000000000",
10387 => "0000000000000000",10388 => "0000000000000000",
10389 => "0000000000000000",10390 => "0000000000000000",
10391 => "0000000000000000",10392 => "0000000000000000",
10393 => "0000000000000000",10394 => "0000000000000000",
10395 => "0000000000000000",10396 => "0000000000000000",
10397 => "0000000000000000",10398 => "0000000000000000",
10399 => "0000000000000000",10400 => "0000000000000000",
10401 => "0000000000000000",10402 => "0000000000000000",
10403 => "0000000000000000",10404 => "0000000000000000",
10405 => "0000000000000000",10406 => "0000000000000000",
10407 => "0000000000000000",10408 => "0000000000000000",
10409 => "0000000000000000",10410 => "0000000000000000",
10411 => "0000000000000000",10412 => "0000000000000000",
10413 => "0000000000000000",10414 => "0000000000000000",
10415 => "0000000000000000",10416 => "0000000000000000",
10417 => "0000000000000000",10418 => "0000000000000000",
10419 => "0000000000000000",10420 => "0000000000000000",
10421 => "0000000000000000",10422 => "0000000000000000",
10423 => "0000000000000000",10424 => "0000000000000000",
10425 => "0000000000000000",10426 => "0000000000000000",
10427 => "0000000000000000",10428 => "0000000000000000",
10429 => "0000000000000000",10430 => "0000000000000000",
10431 => "0000000000000000",10432 => "0000000000000000",
10433 => "0000000000000000",10434 => "0000000000000000",
10435 => "0000000000000000",10436 => "0000000000000000",
10437 => "0000000000000000",10438 => "0000000000000000",
10439 => "0000000000000000",10440 => "0000000000000000",
10441 => "0000000000000000",10442 => "0000000000000000",
10443 => "0000000000000000",10444 => "0000000000000000",
10445 => "0000000000000000",10446 => "0000000000000000",
10447 => "0000000000000000",10448 => "0000000000000000",
10449 => "0000000000000000",10450 => "0000000000000000",
10451 => "0000000000000000",10452 => "0000000000000000",
10453 => "0000000000000000",10454 => "0000000000000000",
10455 => "0000000000000000",10456 => "0000000000000000",
10457 => "0000000000000000",10458 => "0000000000000000",
10459 => "0000000000000000",10460 => "0000000000000000",
10461 => "0000000000000000",10462 => "0000000000000000",
10463 => "0000000000000000",10464 => "0000000000000000",
10465 => "0000000000000000",10466 => "0000000000000000",
10467 => "0000000000000000",10468 => "0000000000000000",
10469 => "0000000000000000",10470 => "0000000000000000",
10471 => "0000000000000000",10472 => "0000000000000000",
10473 => "0000000000000000",10474 => "0000000000000000",
10475 => "0000000000000000",10476 => "0000000000000000",
10477 => "0000000000000000",10478 => "0000000000000000",
10479 => "0000000000000000",10480 => "0000000000000000",
10481 => "0000000000000000",10482 => "0000000000000000",
10483 => "0000000000000000",10484 => "0000000000000000",
10485 => "0000000000000000",10486 => "0000000000000000",
10487 => "0000000000000000",10488 => "0000000000000000",
10489 => "0000000000000000",10490 => "0000000000000000",
10491 => "0000000000000000",10492 => "0000000000000000",
10493 => "0000000000000000",10494 => "0000000000000000",
10495 => "0000000000000000",10496 => "0000000000000000",
10497 => "0000000000000000",10498 => "0000000000000000",
10499 => "0000000000000000",10500 => "0000000000000000",
10501 => "0000000000000000",10502 => "0000000000000000",
10503 => "0000000000000000",10504 => "0000000000000000",
10505 => "0000000000000000",10506 => "0000000000000000",
10507 => "0000000000000000",10508 => "0000000000000000",
10509 => "0000000000000000",10510 => "0000000000000000",
10511 => "0000000000000000",10512 => "0000000000000000",
10513 => "0000000000000000",10514 => "0000000000000000",
10515 => "0000000000000000",10516 => "0000000000000000",
10517 => "0000000000000000",10518 => "0000000000000000",
10519 => "0000000000000000",10520 => "0000000000000000",
10521 => "0000000000000000",10522 => "0000000000000000",
10523 => "0000000000000000",10524 => "0000000000000000",
10525 => "0000000000000000",10526 => "0000000000000000",
10527 => "0000000000000000",10528 => "0000000000000000",
10529 => "0000000000000000",10530 => "0000000000000000",
10531 => "0000000000000000",10532 => "0000000000000000",
10533 => "0000000000000000",10534 => "0000000000000000",
10535 => "0000000000000000",10536 => "0000000000000000",
10537 => "0000000000000000",10538 => "0000000000000000",
10539 => "0000000000000000",10540 => "0000000000000000",
10541 => "0000000000000000",10542 => "0000000000000000",
10543 => "0000000000000000",10544 => "0000000000000000",
10545 => "0000000000000000",10546 => "0000000000000000",
10547 => "0000000000000000",10548 => "0000000000000000",
10549 => "0000000000000000",10550 => "0000000000000000",
10551 => "0000000000000000",10552 => "0000000000000000",
10553 => "0000000000000000",10554 => "0000000000000000",
10555 => "0000000000000000",10556 => "0000000000000000",
10557 => "0000000000000000",10558 => "0000000000000000",
10559 => "0000000000000000",10560 => "0000000000000000",
10561 => "0000000000000000",10562 => "0000000000000000",
10563 => "0000000000000000",10564 => "0000000000000000",
10565 => "0000000000000000",10566 => "0000000000000000",
10567 => "0000000000000000",10568 => "0000000000000000",
10569 => "0000000000000000",10570 => "0000000000000000",
10571 => "0000000000000000",10572 => "0000000000000000",
10573 => "0000000000000000",10574 => "0000000000000000",
10575 => "0000000000000000",10576 => "0000000000000000",
10577 => "0000000000000000",10578 => "0000000000000000",
10579 => "0000000000000000",10580 => "0000000000000000",
10581 => "0000000000000000",10582 => "0000000000000000",
10583 => "0000000000000000",10584 => "0000000000000000",
10585 => "0000000000000000",10586 => "0000000000000000",
10587 => "0000000000000000",10588 => "0000000000000000",
10589 => "0000000000000000",10590 => "0000000000000000",
10591 => "0000000000000000",10592 => "0000000000000000",
10593 => "0000000000000000",10594 => "0000000000000000",
10595 => "0000000000000000",10596 => "0000000000000000",
10597 => "0000000000000000",10598 => "0000000000000000",
10599 => "0000000000000000",10600 => "0000000000000000",
10601 => "0000000000000000",10602 => "0000000000000000",
10603 => "0000000000000000",10604 => "0000000000000000",
10605 => "0000000000000000",10606 => "0000000000000000",
10607 => "0000000000000000",10608 => "0000000000000000",
10609 => "0000000000000000",10610 => "0000000000000000",
10611 => "0000000000000000",10612 => "0000000000000000",
10613 => "0000000000000000",10614 => "0000000000000000",
10615 => "0000000000000000",10616 => "0000000000000000",
10617 => "0000000000000000",10618 => "0000000000000000",
10619 => "0000000000000000",10620 => "0000000000000000",
10621 => "0000000000000000",10622 => "0000000000000000",
10623 => "0000000000000000",10624 => "0000000000000000",
10625 => "0000000000000000",10626 => "0000000000000000",
10627 => "0000000000000000",10628 => "0000000000000000",
10629 => "0000000000000000",10630 => "0000000000000000",
10631 => "0000000000000000",10632 => "0000000000000000",
10633 => "0000000000000000",10634 => "0000000000000000",
10635 => "0000000000000000",10636 => "0000000000000000",
10637 => "0000000000000000",10638 => "0000000000000000",
10639 => "0000000000000000",10640 => "0000000000000000",
10641 => "0000000000000000",10642 => "0000000000000000",
10643 => "0000000000000000",10644 => "0000000000000000",
10645 => "0000000000000000",10646 => "0000000000000000",
10647 => "0000000000000000",10648 => "0000000000000000",
10649 => "0000000000000000",10650 => "0000000000000000",
10651 => "0000000000000000",10652 => "0000000000000000",
10653 => "0000000000000000",10654 => "0000000000000000",
10655 => "0000000000000000",10656 => "0000000000000000",
10657 => "0000000000000000",10658 => "0000000000000000",
10659 => "0000000000000000",10660 => "0000000000000000",
10661 => "0000000000000000",10662 => "0000000000000000",
10663 => "0000000000000000",10664 => "0000000000000000",
10665 => "0000000000000000",10666 => "0000000000000000",
10667 => "0000000000000000",10668 => "0000000000000000",
10669 => "0000000000000000",10670 => "0000000000000000",
10671 => "0000000000000000",10672 => "0000000000000000",
10673 => "0000000000000000",10674 => "0000000000000000",
10675 => "0000000000000000",10676 => "0000000000000000",
10677 => "0000000000000000",10678 => "0000000000000000",
10679 => "0000000000000000",10680 => "0000000000000000",
10681 => "0000000000000000",10682 => "0000000000000000",
10683 => "0000000000000000",10684 => "0000000000000000",
10685 => "0000000000000000",10686 => "0000000000000000",
10687 => "0000000000000000",10688 => "0000000000000000",
10689 => "0000000000000000",10690 => "0000000000000000",
10691 => "0000000000000000",10692 => "0000000000000000",
10693 => "0000000000000000",10694 => "0000000000000000",
10695 => "0000000000000000",10696 => "0000000000000000",
10697 => "0000000000000000",10698 => "0000000000000000",
10699 => "0000000000000000",10700 => "0000000000000000",
10701 => "0000000000000000",10702 => "0000000000000000",
10703 => "0000000000000000",10704 => "0000000000000000",
10705 => "0000000000000000",10706 => "0000000000000000",
10707 => "0000000000000000",10708 => "0000000000000000",
10709 => "0000000000000000",10710 => "0000000000000000",
10711 => "0000000000000000",10712 => "0000000000000000",
10713 => "0000000000000000",10714 => "0000000000000000",
10715 => "0000000000000000",10716 => "0000000000000000",
10717 => "0000000000000000",10718 => "0000000000000000",
10719 => "0000000000000000",10720 => "0000000000000000",
10721 => "0000000000000000",10722 => "0000000000000000",
10723 => "0000000000000000",10724 => "0000000000000000",
10725 => "0000000000000000",10726 => "0000000000000000",
10727 => "0000000000000000",10728 => "0000000000000000",
10729 => "0000000000000000",10730 => "0000000000000000",
10731 => "0000000000000000",10732 => "0000000000000000",
10733 => "0000000000000000",10734 => "0000000000000000",
10735 => "0000000000000000",10736 => "0000000000000000",
10737 => "0000000000000000",10738 => "0000000000000000",
10739 => "0000000000000000",10740 => "0000000000000000",
10741 => "0000000000000000",10742 => "0000000000000000",
10743 => "0000000000000000",10744 => "0000000000000000",
10745 => "0000000000000000",10746 => "0000000000000000",
10747 => "0000000000000000",10748 => "0000000000000000",
10749 => "0000000000000000",10750 => "0000000000000000",
10751 => "0000000000000000",10752 => "0000000000000000",
10753 => "0000000000000000",10754 => "0000000000000000",
10755 => "0000000000000000",10756 => "0000000000000000",
10757 => "0000000000000000",10758 => "0000000000000000",
10759 => "0000000000000000",10760 => "0000000000000000",
10761 => "0000000000000000",10762 => "0000000000000000",
10763 => "0000000000000000",10764 => "0000000000000000",
10765 => "0000000000000000",10766 => "0000000000000000",
10767 => "0000000000000000",10768 => "0000000000000000",
10769 => "0000000000000000",10770 => "0000000000000000",
10771 => "0000000000000000",10772 => "0000000000000000",
10773 => "0000000000000000",10774 => "0000000000000000",
10775 => "0000000000000000",10776 => "0000000000000000",
10777 => "0000000000000000",10778 => "0000000000000000",
10779 => "0000000000000000",10780 => "0000000000000000",
10781 => "0000000000000000",10782 => "0000000000000000",
10783 => "0000000000000000",10784 => "0000000000000000",
10785 => "0000000000000000",10786 => "0000000000000000",
10787 => "0000000000000000",10788 => "0000000000000000",
10789 => "0000000000000000",10790 => "0000000000000000",
10791 => "0000000000000000",10792 => "0000000000000000",
10793 => "0000000000000000",10794 => "0000000000000000",
10795 => "0000000000000000",10796 => "0000000000000000",
10797 => "0000000000000000",10798 => "0000000000000000",
10799 => "0000000000000000",10800 => "0000000000000000",
10801 => "0000000000000000",10802 => "0000000000000000",
10803 => "0000000000000000",10804 => "0000000000000000",
10805 => "0000000000000000",10806 => "0000000000000000",
10807 => "0000000000000000",10808 => "0000000000000000",
10809 => "0000000000000000",10810 => "0000000000000000",
10811 => "0000000000000000",10812 => "0000000000000000",
10813 => "0000000000000000",10814 => "0000000000000000",
10815 => "0000000000000000",10816 => "0000000000000000",
10817 => "0000000000000000",10818 => "0000000000000000",
10819 => "0000000000000000",10820 => "0000000000000000",
10821 => "0000000000000000",10822 => "0000000000000000",
10823 => "0000000000000000",10824 => "0000000000000000",
10825 => "0000000000000000",10826 => "0000000000000000",
10827 => "0000000000000000",10828 => "0000000000000000",
10829 => "0000000000000000",10830 => "0000000000000000",
10831 => "0000000000000000",10832 => "0000000000000000",
10833 => "0000000000000000",10834 => "0000000000000000",
10835 => "0000000000000000",10836 => "0000000000000000",
10837 => "0000000000000000",10838 => "0000000000000000",
10839 => "0000000000000000",10840 => "0000000000000000",
10841 => "0000000000000000",10842 => "0000000000000000",
10843 => "0000000000000000",10844 => "0000000000000000",
10845 => "0000000000000000",10846 => "0000000000000000",
10847 => "0000000000000000",10848 => "0000000000000000",
10849 => "0000000000000000",10850 => "0000000000000000",
10851 => "0000000000000000",10852 => "0000000000000000",
10853 => "0000000000000000",10854 => "0000000000000000",
10855 => "0000000000000000",10856 => "0000000000000000",
10857 => "0000000000000000",10858 => "0000000000000000",
10859 => "0000000000000000",10860 => "0000000000000000",
10861 => "0000000000000000",10862 => "0000000000000000",
10863 => "0000000000000000",10864 => "0000000000000000",
10865 => "0000000000000000",10866 => "0000000000000000",
10867 => "0000000000000000",10868 => "0000000000000000",
10869 => "0000000000000000",10870 => "0000000000000000",
10871 => "0000000000000000",10872 => "0000000000000000",
10873 => "0000000000000000",10874 => "0000000000000000",
10875 => "0000000000000000",10876 => "0000000000000000",
10877 => "0000000000000000",10878 => "0000000000000000",
10879 => "0000000000000000",10880 => "0000000000000000",
10881 => "0000000000000000",10882 => "0000000000000000",
10883 => "0000000000000000",10884 => "0000000000000000",
10885 => "0000000000000000",10886 => "0000000000000000",
10887 => "0000000000000000",10888 => "0000000000000000",
10889 => "0000000000000000",10890 => "0000000000000000",
10891 => "0000000000000000",10892 => "0000000000000000",
10893 => "0000000000000000",10894 => "0000000000000000",
10895 => "0000000000000000",10896 => "0000000000000000",
10897 => "0000000000000000",10898 => "0000000000000000",
10899 => "0000000000000000",10900 => "0000000000000000",
10901 => "0000000000000000",10902 => "0000000000000000",
10903 => "0000000000000000",10904 => "0000000000000000",
10905 => "0000000000000000",10906 => "0000000000000000",
10907 => "0000000000000000",10908 => "0000000000000000",
10909 => "0000000000000000",10910 => "0000000000000000",
10911 => "0000000000000000",10912 => "0000000000000000",
10913 => "0000000000000000",10914 => "0000000000000000",
10915 => "0000000000000000",10916 => "0000000000000000",
10917 => "0000000000000000",10918 => "0000000000000000",
10919 => "0000000000000000",10920 => "0000000000000000",
10921 => "0000000000000000",10922 => "0000000000000000",
10923 => "0000000000000000",10924 => "0000000000000000",
10925 => "0000000000000000",10926 => "0000000000000000",
10927 => "0000000000000000",10928 => "0000000000000000",
10929 => "0000000000000000",10930 => "0000000000000000",
10931 => "0000000000000000",10932 => "0000000000000000",
10933 => "0000000000000000",10934 => "0000000000000000",
10935 => "0000000000000000",10936 => "0000000000000000",
10937 => "0000000000000000",10938 => "0000000000000000",
10939 => "0000000000000000",10940 => "0000000000000000",
10941 => "0000000000000000",10942 => "0000000000000000",
10943 => "0000000000000000",10944 => "0000000000000000",
10945 => "0000000000000000",10946 => "0000000000000000",
10947 => "0000000000000000",10948 => "0000000000000000",
10949 => "0000000000000000",10950 => "0000000000000000",
10951 => "0000000000000000",10952 => "0000000000000000",
10953 => "0000000000000000",10954 => "0000000000000000",
10955 => "0000000000000000",10956 => "0000000000000000",
10957 => "0000000000000000",10958 => "0000000000000000",
10959 => "0000000000000000",10960 => "0000000000000000",
10961 => "0000000000000000",10962 => "0000000000000000",
10963 => "0000000000000000",10964 => "0000000000000000",
10965 => "0000000000000000",10966 => "0000000000000000",
10967 => "0000000000000000",10968 => "0000000000000000",
10969 => "0000000000000000",10970 => "0000000000000000",
10971 => "0000000000000000",10972 => "0000000000000000",
10973 => "0000000000000000",10974 => "0000000000000000",
10975 => "0000000000000000",10976 => "0000000000000000",
10977 => "0000000000000000",10978 => "0000000000000000",
10979 => "0000000000000000",10980 => "0000000000000000",
10981 => "0000000000000000",10982 => "0000000000000000",
10983 => "0000000000000000",10984 => "0000000000000000",
10985 => "0000000000000000",10986 => "0000000000000000",
10987 => "0000000000000000",10988 => "0000000000000000",
10989 => "0000000000000000",10990 => "0000000000000000",
10991 => "0000000000000000",10992 => "0000000000000000",
10993 => "0000000000000000",10994 => "0000000000000000",
10995 => "0000000000000000",10996 => "0000000000000000",
10997 => "0000000000000000",10998 => "0000000000000000",
10999 => "0000000000000000",11000 => "0000000000000000",
11001 => "0000000000000000",11002 => "0000000000000000",
11003 => "0000000000000000",11004 => "0000000000000000",
11005 => "0000000000000000",11006 => "0000000000000000",
11007 => "0000000000000000",11008 => "0000000000000000",
11009 => "0000000000000000",11010 => "0000000000000000",
11011 => "0000000000000000",11012 => "0000000000000000",
11013 => "0000000000000000",11014 => "0000000000000000",
11015 => "0000000000000000",11016 => "0000000000000000",
11017 => "0000000000000000",11018 => "0000000000000000",
11019 => "0000000000000000",11020 => "0000000000000000",
11021 => "0000000000000000",11022 => "0000000000000000",
11023 => "0000000000000000",11024 => "0000000000000000",
11025 => "0000000000000000",11026 => "0000000000000000",
11027 => "0000000000000000",11028 => "0000000000000000",
11029 => "0000000000000000",11030 => "0000000000000000",
11031 => "0000000000000000",11032 => "0000000000000000",
11033 => "0000000000000000",11034 => "0000000000000000",
11035 => "0000000000000000",11036 => "0000000000000000",
11037 => "0000000000000000",11038 => "0000000000000000",
11039 => "0000000000000000",11040 => "0000000000000000",
11041 => "0000000000000000",11042 => "0000000000000000",
11043 => "0000000000000000",11044 => "0000000000000000",
11045 => "0000000000000000",11046 => "0000000000000000",
11047 => "0000000000000000",11048 => "0000000000000000",
11049 => "0000000000000000",11050 => "0000000000000000",
11051 => "0000000000000000",11052 => "0000000000000000",
11053 => "0000000000000000",11054 => "0000000000000000",
11055 => "0000000000000000",11056 => "0000000000000000",
11057 => "0000000000000000",11058 => "0000000000000000",
11059 => "0000000000000000",11060 => "0000000000000000",
11061 => "0000000000000000",11062 => "0000000000000000",
11063 => "0000000000000000",11064 => "0000000000000000",
11065 => "0000000000000000",11066 => "0000000000000000",
11067 => "0000000000000000",11068 => "0000000000000000",
11069 => "0000000000000000",11070 => "0000000000000000",
11071 => "0000000000000000",11072 => "0000000000000000",
11073 => "0000000000000000",11074 => "0000000000000000",
11075 => "0000000000000000",11076 => "0000000000000000",
11077 => "0000000000000000",11078 => "0000000000000000",
11079 => "0000000000000000",11080 => "0000000000000000",
11081 => "0000000000000000",11082 => "0000000000000000",
11083 => "0000000000000000",11084 => "0000000000000000",
11085 => "0000000000000000",11086 => "0000000000000000",
11087 => "0000000000000000",11088 => "0000000000000000",
11089 => "0000000000000000",11090 => "0000000000000000",
11091 => "0000000000000000",11092 => "0000000000000000",
11093 => "0000000000000000",11094 => "0000000000000000",
11095 => "0000000000000000",11096 => "0000000000000000",
11097 => "0000000000000000",11098 => "0000000000000000",
11099 => "0000000000000000",11100 => "0000000000000000",
11101 => "0000000000000000",11102 => "0000000000000000",
11103 => "0000000000000000",11104 => "0000000000000000",
11105 => "0000000000000000",11106 => "0000000000000000",
11107 => "0000000000000000",11108 => "0000000000000000",
11109 => "0000000000000000",11110 => "0000000000000000",
11111 => "0000000000000000",11112 => "0000000000000000",
11113 => "0000000000000000",11114 => "0000000000000000",
11115 => "0000000000000000",11116 => "0000000000000000",
11117 => "0000000000000000",11118 => "0000000000000000",
11119 => "0000000000000000",11120 => "0000000000000000",
11121 => "0000000000000000",11122 => "0000000000000000",
11123 => "0000000000000000",11124 => "0000000000000000",
11125 => "0000000000000000",11126 => "0000000000000000",
11127 => "0000000000000000",11128 => "0000000000000000",
11129 => "0000000000000000",11130 => "0000000000000000",
11131 => "0000000000000000",11132 => "0000000000000000",
11133 => "0000000000000000",11134 => "0000000000000000",
11135 => "0000000000000000",11136 => "0000000000000000",
11137 => "0000000000000000",11138 => "0000000000000000",
11139 => "0000000000000000",11140 => "0000000000000000",
11141 => "0000000000000000",11142 => "0000000000000000",
11143 => "0000000000000000",11144 => "0000000000000000",
11145 => "0000000000000000",11146 => "0000000000000000",
11147 => "0000000000000000",11148 => "0000000000000000",
11149 => "0000000000000000",11150 => "0000000000000000",
11151 => "0000000000000000",11152 => "0000000000000000",
11153 => "0000000000000000",11154 => "0000000000000000",
11155 => "0000000000000000",11156 => "0000000000000000",
11157 => "0000000000000000",11158 => "0000000000000000",
11159 => "0000000000000000",11160 => "0000000000000000",
11161 => "0000000000000000",11162 => "0000000000000000",
11163 => "0000000000000000",11164 => "0000000000000000",
11165 => "0000000000000000",11166 => "0000000000000000",
11167 => "0000000000000000",11168 => "0000000000000000",
11169 => "0000000000000000",11170 => "0000000000000000",
11171 => "0000000000000000",11172 => "0000000000000000",
11173 => "0000000000000000",11174 => "0000000000000000",
11175 => "0000000000000000",11176 => "0000000000000000",
11177 => "0000000000000000",11178 => "0000000000000000",
11179 => "0000000000000000",11180 => "0000000000000000",
11181 => "0000000000000000",11182 => "0000000000000000",
11183 => "0000000000000000",11184 => "0000000000000000",
11185 => "0000000000000000",11186 => "0000000000000000",
11187 => "0000000000000000",11188 => "0000000000000000",
11189 => "0000000000000000",11190 => "0000000000000000",
11191 => "0000000000000000",11192 => "0000000000000000",
11193 => "0000000000000000",11194 => "0000000000000000",
11195 => "0000000000000000",11196 => "0000000000000000",
11197 => "0000000000000000",11198 => "0000000000000000",
11199 => "0000000000000000",11200 => "0000000000000000",
11201 => "0000000000000000",11202 => "0000000000000000",
11203 => "0000000000000000",11204 => "0000000000000000",
11205 => "0000000000000000",11206 => "0000000000000000",
11207 => "0000000000000000",11208 => "0000000000000000",
11209 => "0000000000000000",11210 => "0000000000000000",
11211 => "0000000000000000",11212 => "0000000000000000",
11213 => "0000000000000000",11214 => "0000000000000000",
11215 => "0000000000000000",11216 => "0000000000000000",
11217 => "0000000000000000",11218 => "0000000000000000",
11219 => "0000000000000000",11220 => "0000000000000000",
11221 => "0000000000000000",11222 => "0000000000000000",
11223 => "0000000000000000",11224 => "0000000000000000",
11225 => "0000000000000000",11226 => "0000000000000000",
11227 => "0000000000000000",11228 => "0000000000000000",
11229 => "0000000000000000",11230 => "0000000000000000",
11231 => "0000000000000000",11232 => "0000000000000000",
11233 => "0000000000000000",11234 => "0000000000000000",
11235 => "0000000000000000",11236 => "0000000000000000",
11237 => "0000000000000000",11238 => "0000000000000000",
11239 => "0000000000000000",11240 => "0000000000000000",
11241 => "0000000000000000",11242 => "0000000000000000",
11243 => "0000000000000000",11244 => "0000000000000000",
11245 => "0000000000000000",11246 => "0000000000000000",
11247 => "0000000000000000",11248 => "0000000000000000",
11249 => "0000000000000000",11250 => "0000000000000000",
11251 => "0000000000000000",11252 => "0000000000000000",
11253 => "0000000000000000",11254 => "0000000000000000",
11255 => "0000000000000000",11256 => "0000000000000000",
11257 => "0000000000000000",11258 => "0000000000000000",
11259 => "0000000000000000",11260 => "0000000000000000",
11261 => "0000000000000000",11262 => "0000000000000000",
11263 => "0000000000000000",11264 => "0000000000000000",
11265 => "0000000000000000",11266 => "0000000000000000",
11267 => "0000000000000000",11268 => "0000000000000000",
11269 => "0000000000000000",11270 => "0000000000000000",
11271 => "0000000000000000",11272 => "0000000000000000",
11273 => "0000000000000000",11274 => "0000000000000000",
11275 => "0000000000000000",11276 => "0000000000000000",
11277 => "0000000000000000",11278 => "0000000000000000",
11279 => "0000000000000000",11280 => "0000000000000000",
11281 => "0000000000000000",11282 => "0000000000000000",
11283 => "0000000000000000",11284 => "0000000000000000",
11285 => "0000000000000000",11286 => "0000000000000000",
11287 => "0000000000000000",11288 => "0000000000000000",
11289 => "0000000000000000",11290 => "0000000000000000",
11291 => "0000000000000000",11292 => "0000000000000000",
11293 => "0000000000000000",11294 => "0000000000000000",
11295 => "0000000000000000",11296 => "0000000000000000",
11297 => "0000000000000000",11298 => "0000000000000000",
11299 => "0000000000000000",11300 => "0000000000000000",
11301 => "0000000000000000",11302 => "0000000000000000",
11303 => "0000000000000000",11304 => "0000000000000000",
11305 => "0000000000000000",11306 => "0000000000000000",
11307 => "0000000000000000",11308 => "0000000000000000",
11309 => "0000000000000000",11310 => "0000000000000000",
11311 => "0000000000000000",11312 => "0000000000000000",
11313 => "0000000000000000",11314 => "0000000000000000",
11315 => "0000000000000000",11316 => "0000000000000000",
11317 => "0000000000000000",11318 => "0000000000000000",
11319 => "0000000000000000",11320 => "0000000000000000",
11321 => "0000000000000000",11322 => "0000000000000000",
11323 => "0000000000000000",11324 => "0000000000000000",
11325 => "0000000000000000",11326 => "0000000000000000",
11327 => "0000000000000000",11328 => "0000000000000000",
11329 => "0000000000000000",11330 => "0000000000000000",
11331 => "0000000000000000",11332 => "0000000000000000",
11333 => "0000000000000000",11334 => "0000000000000000",
11335 => "0000000000000000",11336 => "0000000000000000",
11337 => "0000000000000000",11338 => "0000000000000000",
11339 => "0000000000000000",11340 => "0000000000000000",
11341 => "0000000000000000",11342 => "0000000000000000",
11343 => "0000000000000000",11344 => "0000000000000000",
11345 => "0000000000000000",11346 => "0000000000000000",
11347 => "0000000000000000",11348 => "0000000000000000",
11349 => "0000000000000000",11350 => "0000000000000000",
11351 => "0000000000000000",11352 => "0000000000000000",
11353 => "0000000000000000",11354 => "0000000000000000",
11355 => "0000000000000000",11356 => "0000000000000000",
11357 => "0000000000000000",11358 => "0000000000000000",
11359 => "0000000000000000",11360 => "0000000000000000",
11361 => "0000000000000000",11362 => "0000000000000000",
11363 => "0000000000000000",11364 => "0000000000000000",
11365 => "0000000000000000",11366 => "0000000000000000",
11367 => "0000000000000000",11368 => "0000000000000000",
11369 => "0000000000000000",11370 => "0000000000000000",
11371 => "0000000000000000",11372 => "0000000000000000",
11373 => "0000000000000000",11374 => "0000000000000000",
11375 => "0000000000000000",11376 => "0000000000000000",
11377 => "0000000000000000",11378 => "0000000000000000",
11379 => "0000000000000000",11380 => "0000000000000000",
11381 => "0000000000000000",11382 => "0000000000000000",
11383 => "0000000000000000",11384 => "0000000000000000",
11385 => "0000000000000000",11386 => "0000000000000000",
11387 => "0000000000000000",11388 => "0000000000000000",
11389 => "0000000000000000",11390 => "0000000000000000",
11391 => "0000000000000000",11392 => "0000000000000000",
11393 => "0000000000000000",11394 => "0000000000000000",
11395 => "0000000000000000",11396 => "0000000000000000",
11397 => "0000000000000000",11398 => "0000000000000000",
11399 => "0000000000000000",11400 => "0000000000000000",
11401 => "0000000000000000",11402 => "0000000000000000",
11403 => "0000000000000000",11404 => "0000000000000000",
11405 => "0000000000000000",11406 => "0000000000000000",
11407 => "0000000000000000",11408 => "0000000000000000",
11409 => "0000000000000000",11410 => "0000000000000000",
11411 => "0000000000000000",11412 => "0000000000000000",
11413 => "0000000000000000",11414 => "0000000000000000",
11415 => "0000000000000000",11416 => "0000000000000000",
11417 => "0000000000000000",11418 => "0000000000000000",
11419 => "0000000000000000",11420 => "0000000000000000",
11421 => "0000000000000000",11422 => "0000000000000000",
11423 => "0000000000000000",11424 => "0000000000000000",
11425 => "0000000000000000",11426 => "0000000000000000",
11427 => "0000000000000000",11428 => "0000000000000000",
11429 => "0000000000000000",11430 => "0000000000000000",
11431 => "0000000000000000",11432 => "0000000000000000",
11433 => "0000000000000000",11434 => "0000000000000000",
11435 => "0000000000000000",11436 => "0000000000000000",
11437 => "0000000000000000",11438 => "0000000000000000",
11439 => "0000000000000000",11440 => "0000000000000000",
11441 => "0000000000000000",11442 => "0000000000000000",
11443 => "0000000000000000",11444 => "0000000000000000",
11445 => "0000000000000000",11446 => "0000000000000000",
11447 => "0000000000000000",11448 => "0000000000000000",
11449 => "0000000000000000",11450 => "0000000000000000",
11451 => "0000000000000000",11452 => "0000000000000000",
11453 => "0000000000000000",11454 => "0000000000000000",
11455 => "0000000000000000",11456 => "0000000000000000",
11457 => "0000000000000000",11458 => "0000000000000000",
11459 => "0000000000000000",11460 => "0000000000000000",
11461 => "0000000000000000",11462 => "0000000000000000",
11463 => "0000000000000000",11464 => "0000000000000000",
11465 => "0000000000000000",11466 => "0000000000000000",
11467 => "0000000000000000",11468 => "0000000000000000",
11469 => "0000000000000000",11470 => "0000000000000000",
11471 => "0000000000000000",11472 => "0000000000000000",
11473 => "0000000000000000",11474 => "0000000000000000",
11475 => "0000000000000000",11476 => "0000000000000000",
11477 => "0000000000000000",11478 => "0000000000000000",
11479 => "0000000000000000",11480 => "0000000000000000",
11481 => "0000000000000000",11482 => "0000000000000000",
11483 => "0000000000000000",11484 => "0000000000000000",
11485 => "0000000000000000",11486 => "0000000000000000",
11487 => "0000000000000000",11488 => "0000000000000000",
11489 => "0000000000000000",11490 => "0000000000000000",
11491 => "0000000000000000",11492 => "0000000000000000",
11493 => "0000000000000000",11494 => "0000000000000000",
11495 => "0000000000000000",11496 => "0000000000000000",
11497 => "0000000000000000",11498 => "0000000000000000",
11499 => "0000000000000000",11500 => "0000000000000000",
11501 => "0000000000000000",11502 => "0000000000000000",
11503 => "0000000000000000",11504 => "0000000000000000",
11505 => "0000000000000000",11506 => "0000000000000000",
11507 => "0000000000000000",11508 => "0000000000000000",
11509 => "0000000000000000",11510 => "0000000000000000",
11511 => "0000000000000000",11512 => "0000000000000000",
11513 => "0000000000000000",11514 => "0000000000000000",
11515 => "0000000000000000",11516 => "0000000000000000",
11517 => "0000000000000000",11518 => "0000000000000000",
11519 => "0000000000000000",11520 => "0000000000000000",
11521 => "0000000000000000",11522 => "0000000000000000",
11523 => "0000000000000000",11524 => "0000000000000000",
11525 => "0000000000000000",11526 => "0000000000000000",
11527 => "0000000000000000",11528 => "0000000000000000",
11529 => "0000000000000000",11530 => "0000000000000000",
11531 => "0000000000000000",11532 => "0000000000000000",
11533 => "0000000000000000",11534 => "0000000000000000",
11535 => "0000000000000000",11536 => "0000000000000000",
11537 => "0000000000000000",11538 => "0000000000000000",
11539 => "0000000000000000",11540 => "0000000000000000",
11541 => "0000000000000000",11542 => "0000000000000000",
11543 => "0000000000000000",11544 => "0000000000000000",
11545 => "0000000000000000",11546 => "0000000000000000",
11547 => "0000000000000000",11548 => "0000000000000000",
11549 => "0000000000000000",11550 => "0000000000000000",
11551 => "0000000000000000",11552 => "0000000000000000",
11553 => "0000000000000000",11554 => "0000000000000000",
11555 => "0000000000000000",11556 => "0000000000000000",
11557 => "0000000000000000",11558 => "0000000000000000",
11559 => "0000000000000000",11560 => "0000000000000000",
11561 => "0000000000000000",11562 => "0000000000000000",
11563 => "0000000000000000",11564 => "0000000000000000",
11565 => "0000000000000000",11566 => "0000000000000000",
11567 => "0000000000000000",11568 => "0000000000000000",
11569 => "0000000000000000",11570 => "0000000000000000",
11571 => "0000000000000000",11572 => "0000000000000000",
11573 => "0000000000000000",11574 => "0000000000000000",
11575 => "0000000000000000",11576 => "0000000000000000",
11577 => "0000000000000000",11578 => "0000000000000000",
11579 => "0000000000000000",11580 => "0000000000000000",
11581 => "0000000000000000",11582 => "0000000000000000",
11583 => "0000000000000000",11584 => "0000000000000000",
11585 => "0000000000000000",11586 => "0000000000000000",
11587 => "0000000000000000",11588 => "0000000000000000",
11589 => "0000000000000000",11590 => "0000000000000000",
11591 => "0000000000000000",11592 => "0000000000000000",
11593 => "0000000000000000",11594 => "0000000000000000",
11595 => "0000000000000000",11596 => "0000000000000000",
11597 => "0000000000000000",11598 => "0000000000000000",
11599 => "0000000000000000",11600 => "0000000000000000",
11601 => "0000000000000000",11602 => "0000000000000000",
11603 => "0000000000000000",11604 => "0000000000000000",
11605 => "0000000000000000",11606 => "0000000000000000",
11607 => "0000000000000000",11608 => "0000000000000000",
11609 => "0000000000000000",11610 => "0000000000000000",
11611 => "0000000000000000",11612 => "0000000000000000",
11613 => "0000000000000000",11614 => "0000000000000000",
11615 => "0000000000000000",11616 => "0000000000000000",
11617 => "0000000000000000",11618 => "0000000000000000",
11619 => "0000000000000000",11620 => "0000000000000000",
11621 => "0000000000000000",11622 => "0000000000000000",
11623 => "0000000000000000",11624 => "0000000000000000",
11625 => "0000000000000000",11626 => "0000000000000000",
11627 => "0000000000000000",11628 => "0000000000000000",
11629 => "0000000000000000",11630 => "0000000000000000",
11631 => "0000000000000000",11632 => "0000000000000000",
11633 => "0000000000000000",11634 => "0000000000000000",
11635 => "0000000000000000",11636 => "0000000000000000",
11637 => "0000000000000000",11638 => "0000000000000000",
11639 => "0000000000000000",11640 => "0000000000000000",
11641 => "0000000000000000",11642 => "0000000000000000",
11643 => "0000000000000000",11644 => "0000000000000000",
11645 => "0000000000000000",11646 => "0000000000000000",
11647 => "0000000000000000",11648 => "0000000000000000",
11649 => "0000000000000000",11650 => "0000000000000000",
11651 => "0000000000000000",11652 => "0000000000000000",
11653 => "0000000000000000",11654 => "0000000000000000",
11655 => "0000000000000000",11656 => "0000000000000000",
11657 => "0000000000000000",11658 => "0000000000000000",
11659 => "0000000000000000",11660 => "0000000000000000",
11661 => "0000000000000000",11662 => "0000000000000000",
11663 => "0000000000000000",11664 => "0000000000000000",
11665 => "0000000000000000",11666 => "0000000000000000",
11667 => "0000000000000000",11668 => "0000000000000000",
11669 => "0000000000000000",11670 => "0000000000000000",
11671 => "0000000000000000",11672 => "0000000000000000",
11673 => "0000000000000000",11674 => "0000000000000000",
11675 => "0000000000000000",11676 => "0000000000000000",
11677 => "0000000000000000",11678 => "0000000000000000",
11679 => "0000000000000000",11680 => "0000000000000000",
11681 => "0000000000000000",11682 => "0000000000000000",
11683 => "0000000000000000",11684 => "0000000000000000",
11685 => "0000000000000000",11686 => "0000000000000000",
11687 => "0000000000000000",11688 => "0000000000000000",
11689 => "0000000000000000",11690 => "0000000000000000",
11691 => "0000000000000000",11692 => "0000000000000000",
11693 => "0000000000000000",11694 => "0000000000000000",
11695 => "0000000000000000",11696 => "0000000000000000",
11697 => "0000000000000000",11698 => "0000000000000000",
11699 => "0000000000000000",11700 => "0000000000000000",
11701 => "0000000000000000",11702 => "0000000000000000",
11703 => "0000000000000000",11704 => "0000000000000000",
11705 => "0000000000000000",11706 => "0000000000000000",
11707 => "0000000000000000",11708 => "0000000000000000",
11709 => "0000000000000000",11710 => "0000000000000000",
11711 => "0000000000000000",11712 => "0000000000000000",
11713 => "0000000000000000",11714 => "0000000000000000",
11715 => "0000000000000000",11716 => "0000000000000000",
11717 => "0000000000000000",11718 => "0000000000000000",
11719 => "0000000000000000",11720 => "0000000000000000",
11721 => "0000000000000000",11722 => "0000000000000000",
11723 => "0000000000000000",11724 => "0000000000000000",
11725 => "0000000000000000",11726 => "0000000000000000",
11727 => "0000000000000000",11728 => "0000000000000000",
11729 => "0000000000000000",11730 => "0000000000000000",
11731 => "0000000000000000",11732 => "0000000000000000",
11733 => "0000000000000000",11734 => "0000000000000000",
11735 => "0000000000000000",11736 => "0000000000000000",
11737 => "0000000000000000",11738 => "0000000000000000",
11739 => "0000000000000000",11740 => "0000000000000000",
11741 => "0000000000000000",11742 => "0000000000000000",
11743 => "0000000000000000",11744 => "0000000000000000",
11745 => "0000000000000000",11746 => "0000000000000000",
11747 => "0000000000000000",11748 => "0000000000000000",
11749 => "0000000000000000",11750 => "0000000000000000",
11751 => "0000000000000000",11752 => "0000000000000000",
11753 => "0000000000000000",11754 => "0000000000000000",
11755 => "0000000000000000",11756 => "0000000000000000",
11757 => "0000000000000000",11758 => "0000000000000000",
11759 => "0000000000000000",11760 => "0000000000000000",
11761 => "0000000000000000",11762 => "0000000000000000",
11763 => "0000000000000000",11764 => "0000000000000000",
11765 => "0000000000000000",11766 => "0000000000000000",
11767 => "0000000000000000",11768 => "0000000000000000",
11769 => "0000000000000000",11770 => "0000000000000000",
11771 => "0000000000000000",11772 => "0000000000000000",
11773 => "0000000000000000",11774 => "0000000000000000",
11775 => "0000000000000000",11776 => "0000000000000000",
11777 => "0000000000000000",11778 => "0000000000000000",
11779 => "0000000000000000",11780 => "0000000000000000",
11781 => "0000000000000000",11782 => "0000000000000000",
11783 => "0000000000000000",11784 => "0000000000000000",
11785 => "0000000000000000",11786 => "0000000000000000",
11787 => "0000000000000000",11788 => "0000000000000000",
11789 => "0000000000000000",11790 => "0000000000000000",
11791 => "0000000000000000",11792 => "0000000000000000",
11793 => "0000000000000000",11794 => "0000000000000000",
11795 => "0000000000000000",11796 => "0000000000000000",
11797 => "0000000000000000",11798 => "0000000000000000",
11799 => "0000000000000000",11800 => "0000000000000000",
11801 => "0000000000000000",11802 => "0000000000000000",
11803 => "0000000000000000",11804 => "0000000000000000",
11805 => "0000000000000000",11806 => "0000000000000000",
11807 => "0000000000000000",11808 => "0000000000000000",
11809 => "0000000000000000",11810 => "0000000000000000",
11811 => "0000000000000000",11812 => "0000000000000000",
11813 => "0000000000000000",11814 => "0000000000000000",
11815 => "0000000000000000",11816 => "0000000000000000",
11817 => "0000000000000000",11818 => "0000000000000000",
11819 => "0000000000000000",11820 => "0000000000000000",
11821 => "0000000000000000",11822 => "0000000000000000",
11823 => "0000000000000000",11824 => "0000000000000000",
11825 => "0000000000000000",11826 => "0000000000000000",
11827 => "0000000000000000",11828 => "0000000000000000",
11829 => "0000000000000000",11830 => "0000000000000000",
11831 => "0000000000000000",11832 => "0000000000000000",
11833 => "0000000000000000",11834 => "0000000000000000",
11835 => "0000000000000000",11836 => "0000000000000000",
11837 => "0000000000000000",11838 => "0000000000000000",
11839 => "0000000000000000",11840 => "0000000000000000",
11841 => "0000000000000000",11842 => "0000000000000000",
11843 => "0000000000000000",11844 => "0000000000000000",
11845 => "0000000000000000",11846 => "0000000000000000",
11847 => "0000000000000000",11848 => "0000000000000000",
11849 => "0000000000000000",11850 => "0000000000000000",
11851 => "0000000000000000",11852 => "0000000000000000",
11853 => "0000000000000000",11854 => "0000000000000000",
11855 => "0000000000000000",11856 => "0000000000000000",
11857 => "0000000000000000",11858 => "0000000000000000",
11859 => "0000000000000000",11860 => "0000000000000000",
11861 => "0000000000000000",11862 => "0000000000000000",
11863 => "0000000000000000",11864 => "0000000000000000",
11865 => "0000000000000000",11866 => "0000000000000000",
11867 => "0000000000000000",11868 => "0000000000000000",
11869 => "0000000000000000",11870 => "0000000000000000",
11871 => "0000000000000000",11872 => "0000000000000000",
11873 => "0000000000000000",11874 => "0000000000000000",
11875 => "0000000000000000",11876 => "0000000000000000",
11877 => "0000000000000000",11878 => "0000000000000000",
11879 => "0000000000000000",11880 => "0000000000000000",
11881 => "0000000000000000",11882 => "0000000000000000",
11883 => "0000000000000000",11884 => "0000000000000000",
11885 => "0000000000000000",11886 => "0000000000000000",
11887 => "0000000000000000",11888 => "0000000000000000",
11889 => "0000000000000000",11890 => "0000000000000000",
11891 => "0000000000000000",11892 => "0000000000000000",
11893 => "0000000000000000",11894 => "0000000000000000",
11895 => "0000000000000000",11896 => "0000000000000000",
11897 => "0000000000000000",11898 => "0000000000000000",
11899 => "0000000000000000",11900 => "0000000000000000",
11901 => "0000000000000000",11902 => "0000000000000000",
11903 => "0000000000000000",11904 => "0000000000000000",
11905 => "0000000000000000",11906 => "0000000000000000",
11907 => "0000000000000000",11908 => "0000000000000000",
11909 => "0000000000000000",11910 => "0000000000000000",
11911 => "0000000000000000",11912 => "0000000000000000",
11913 => "0000000000000000",11914 => "0000000000000000",
11915 => "0000000000000000",11916 => "0000000000000000",
11917 => "0000000000000000",11918 => "0000000000000000",
11919 => "0000000000000000",11920 => "0000000000000000",
11921 => "0000000000000000",11922 => "0000000000000000",
11923 => "0000000000000000",11924 => "0000000000000000",
11925 => "0000000000000000",11926 => "0000000000000000",
11927 => "0000000000000000",11928 => "0000000000000000",
11929 => "0000000000000000",11930 => "0000000000000000",
11931 => "0000000000000000",11932 => "0000000000000000",
11933 => "0000000000000000",11934 => "0000000000000000",
11935 => "0000000000000000",11936 => "0000000000000000",
11937 => "0000000000000000",11938 => "0000000000000000",
11939 => "0000000000000000",11940 => "0000000000000000",
11941 => "0000000000000000",11942 => "0000000000000000",
11943 => "0000000000000000",11944 => "0000000000000000",
11945 => "0000000000000000",11946 => "0000000000000000",
11947 => "0000000000000000",11948 => "0000000000000000",
11949 => "0000000000000000",11950 => "0000000000000000",
11951 => "0000000000000000",11952 => "0000000000000000",
11953 => "0000000000000000",11954 => "0000000000000000",
11955 => "0000000000000000",11956 => "0000000000000000",
11957 => "0000000000000000",11958 => "0000000000000000",
11959 => "0000000000000000",11960 => "0000000000000000",
11961 => "0000000000000000",11962 => "0000000000000000",
11963 => "0000000000000000",11964 => "0000000000000000",
11965 => "0000000000000000",11966 => "0000000000000000",
11967 => "0000000000000000",11968 => "0000000000000000",
11969 => "0000000000000000",11970 => "0000000000000000",
11971 => "0000000000000000",11972 => "0000000000000000",
11973 => "0000000000000000",11974 => "0000000000000000",
11975 => "0000000000000000",11976 => "0000000000000000",
11977 => "0000000000000000",11978 => "0000000000000000",
11979 => "0000000000000000",11980 => "0000000000000000",
11981 => "0000000000000000",11982 => "0000000000000000",
11983 => "0000000000000000",11984 => "0000000000000000",
11985 => "0000000000000000",11986 => "0000000000000000",
11987 => "0000000000000000",11988 => "0000000000000000",
11989 => "0000000000000000",11990 => "0000000000000000",
11991 => "0000000000000000",11992 => "0000000000000000",
11993 => "0000000000000000",11994 => "0000000000000000",
11995 => "0000000000000000",11996 => "0000000000000000",
11997 => "0000000000000000",11998 => "0000000000000000",
11999 => "0000000000000000",12000 => "0000000000000000",
12001 => "0000000000000000",12002 => "0000000000000000",
12003 => "0000000000000000",12004 => "0000000000000000",
12005 => "0000000000000000",12006 => "0000000000000000",
12007 => "0000000000000000",12008 => "0000000000000000",
12009 => "0000000000000000",12010 => "0000000000000000",
12011 => "0000000000000000",12012 => "0000000000000000",
12013 => "0000000000000000",12014 => "0000000000000000",
12015 => "0000000000000000",12016 => "0000000000000000",
12017 => "0000000000000000",12018 => "0000000000000000",
12019 => "0000000000000000",12020 => "0000000000000000",
12021 => "0000000000000000",12022 => "0000000000000000",
12023 => "0000000000000000",12024 => "0000000000000000",
12025 => "0000000000000000",12026 => "0000000000000000",
12027 => "0000000000000000",12028 => "0000000000000000",
12029 => "0000000000000000",12030 => "0000000000000000",
12031 => "0000000000000000",12032 => "0000000000000000",
12033 => "0000000000000000",12034 => "0000000000000000",
12035 => "0000000000000000",12036 => "0000000000000000",
12037 => "0000000000000000",12038 => "0000000000000000",
12039 => "0000000000000000",12040 => "0000000000000000",
12041 => "0000000000000000",12042 => "0000000000000000",
12043 => "0000000000000000",12044 => "0000000000000000",
12045 => "0000000000000000",12046 => "0000000000000000",
12047 => "0000000000000000",12048 => "0000000000000000",
12049 => "0000000000000000",12050 => "0000000000000000",
12051 => "0000000000000000",12052 => "0000000000000000",
12053 => "0000000000000000",12054 => "0000000000000000",
12055 => "0000000000000000",12056 => "0000000000000000",
12057 => "0000000000000000",12058 => "0000000000000000",
12059 => "0000000000000000",12060 => "0000000000000000",
12061 => "0000000000000000",12062 => "0000000000000000",
12063 => "0000000000000000",12064 => "0000000000000000",
12065 => "0000000000000000",12066 => "0000000000000000",
12067 => "0000000000000000",12068 => "0000000000000000",
12069 => "0000000000000000",12070 => "0000000000000000",
12071 => "0000000000000000",12072 => "0000000000000000",
12073 => "0000000000000000",12074 => "0000000000000000",
12075 => "0000000000000000",12076 => "0000000000000000",
12077 => "0000000000000000",12078 => "0000000000000000",
12079 => "0000000000000000",12080 => "0000000000000000",
12081 => "0000000000000000",12082 => "0000000000000000",
12083 => "0000000000000000",12084 => "0000000000000000",
12085 => "0000000000000000",12086 => "0000000000000000",
12087 => "0000000000000000",12088 => "0000000000000000",
12089 => "0000000000000000",12090 => "0000000000000000",
12091 => "0000000000000000",12092 => "0000000000000000",
12093 => "0000000000000000",12094 => "0000000000000000",
12095 => "0000000000000000",12096 => "0000000000000000",
12097 => "0000000000000000",12098 => "0000000000000000",
12099 => "0000000000000000",12100 => "0000000000000000",
12101 => "0000000000000000",12102 => "0000000000000000",
12103 => "0000000000000000",12104 => "0000000000000000",
12105 => "0000000000000000",12106 => "0000000000000000",
12107 => "0000000000000000",12108 => "0000000000000000",
12109 => "0000000000000000",12110 => "0000000000000000",
12111 => "0000000000000000",12112 => "0000000000000000",
12113 => "0000000000000000",12114 => "0000000000000000",
12115 => "0000000000000000",12116 => "0000000000000000",
12117 => "0000000000000000",12118 => "0000000000000000",
12119 => "0000000000000000",12120 => "0000000000000000",
12121 => "0000000000000000",12122 => "0000000000000000",
12123 => "0000000000000000",12124 => "0000000000000000",
12125 => "0000000000000000",12126 => "0000000000000000",
12127 => "0000000000000000",12128 => "0000000000000000",
12129 => "0000000000000000",12130 => "0000000000000000",
12131 => "0000000000000000",12132 => "0000000000000000",
12133 => "0000000000000000",12134 => "0000000000000000",
12135 => "0000000000000000",12136 => "0000000000000000",
12137 => "0000000000000000",12138 => "0000000000000000",
12139 => "0000000000000000",12140 => "0000000000000000",
12141 => "0000000000000000",12142 => "0000000000000000",
12143 => "0000000000000000",12144 => "0000000000000000",
12145 => "0000000000000000",12146 => "0000000000000000",
12147 => "0000000000000000",12148 => "0000000000000000",
12149 => "0000000000000000",12150 => "0000000000000000",
12151 => "0000000000000000",12152 => "0000000000000000",
12153 => "0000000000000000",12154 => "0000000000000000",
12155 => "0000000000000000",12156 => "0000000000000000",
12157 => "0000000000000000",12158 => "0000000000000000",
12159 => "0000000000000000",12160 => "0000000000000000",
12161 => "0000000000000000",12162 => "0000000000000000",
12163 => "0000000000000000",12164 => "0000000000000000",
12165 => "0000000000000000",12166 => "0000000000000000",
12167 => "0000000000000000",12168 => "0000000000000000",
12169 => "0000000000000000",12170 => "0000000000000000",
12171 => "0000000000000000",12172 => "0000000000000000",
12173 => "0000000000000000",12174 => "0000000000000000",
12175 => "0000000000000000",12176 => "0000000000000000",
12177 => "0000000000000000",12178 => "0000000000000000",
12179 => "0000000000000000",12180 => "0000000000000000",
12181 => "0000000000000000",12182 => "0000000000000000",
12183 => "0000000000000000",12184 => "0000000000000000",
12185 => "0000000000000000",12186 => "0000000000000000",
12187 => "0000000000000000",12188 => "0000000000000000",
12189 => "0000000000000000",12190 => "0000000000000000",
12191 => "0000000000000000",12192 => "0000000000000000",
12193 => "0000000000000000",12194 => "0000000000000000",
12195 => "0000000000000000",12196 => "0000000000000000",
12197 => "0000000000000000",12198 => "0000000000000000",
12199 => "0000000000000000",12200 => "0000000000000000",
12201 => "0000000000000000",12202 => "0000000000000000",
12203 => "0000000000000000",12204 => "0000000000000000",
12205 => "0000000000000000",12206 => "0000000000000000",
12207 => "0000000000000000",12208 => "0000000000000000",
12209 => "0000000000000000",12210 => "0000000000000000",
12211 => "0000000000000000",12212 => "0000000000000000",
12213 => "0000000000000000",12214 => "0000000000000000",
12215 => "0000000000000000",12216 => "0000000000000000",
12217 => "0000000000000000",12218 => "0000000000000000",
12219 => "0000000000000000",12220 => "0000000000000000",
12221 => "0000000000000000",12222 => "0000000000000000",
12223 => "0000000000000000",12224 => "0000000000000000",
12225 => "0000000000000000",12226 => "0000000000000000",
12227 => "0000000000000000",12228 => "0000000000000000",
12229 => "0000000000000000",12230 => "0000000000000000",
12231 => "0000000000000000",12232 => "0000000000000000",
12233 => "0000000000000000",12234 => "0000000000000000",
12235 => "0000000000000000",12236 => "0000000000000000",
12237 => "0000000000000000",12238 => "0000000000000000",
12239 => "0000000000000000",12240 => "0000000000000000",
12241 => "0000000000000000",12242 => "0000000000000000",
12243 => "0000000000000000",12244 => "0000000000000000",
12245 => "0000000000000000",12246 => "0000000000000000",
12247 => "0000000000000000",12248 => "0000000000000000",
12249 => "0000000000000000",12250 => "0000000000000000",
12251 => "0000000000000000",12252 => "0000000000000000",
12253 => "0000000000000000",12254 => "0000000000000000",
12255 => "0000000000000000",12256 => "0000000000000000",
12257 => "0000000000000000",12258 => "0000000000000000",
12259 => "0000000000000000",12260 => "0000000000000000",
12261 => "0000000000000000",12262 => "0000000000000000",
12263 => "0000000000000000",12264 => "0000000000000000",
12265 => "0000000000000000",12266 => "0000000000000000",
12267 => "0000000000000000",12268 => "0000000000000000",
12269 => "0000000000000000",12270 => "0000000000000000",
12271 => "0000000000000000",12272 => "0000000000000000",
12273 => "0000000000000000",12274 => "0000000000000000",
12275 => "0000000000000000",12276 => "0000000000000000",
12277 => "0000000000000000",12278 => "0000000000000000",
12279 => "0000000000000000",12280 => "0000000000000000",
12281 => "0000000000000000",12282 => "0000000000000000",
12283 => "0000000000000000",12284 => "0000000000000000",
12285 => "0000000000000000",12286 => "0000000000000000",
12287 => "0000000000000000",12288 => "0000000000000000",
12289 => "0000000000000000",12290 => "0000000000000000",
12291 => "0000000000000000",12292 => "0000000000000000",
12293 => "0000000000000000",12294 => "0000000000000000",
12295 => "0000000000000000",12296 => "0000000000000000",
12297 => "0000000000000000",12298 => "0000000000000000",
12299 => "0000000000000000",12300 => "0000000000000000",
12301 => "0000000000000000",12302 => "0000000000000000",
12303 => "0000000000000000",12304 => "0000000000000000",
12305 => "0000000000000000",12306 => "0000000000000000",
12307 => "0000000000000000",12308 => "0000000000000000",
12309 => "0000000000000000",12310 => "0000000000000000",
12311 => "0000000000000000",12312 => "0000000000000000",
12313 => "0000000000000000",12314 => "0000000000000000",
12315 => "0000000000000000",12316 => "0000000000000000",
12317 => "0000000000000000",12318 => "0000000000000000",
12319 => "0000000000000000",12320 => "0000000000000000",
12321 => "0000000000000000",12322 => "0000000000000000",
12323 => "0000000000000000",12324 => "0000000000000000",
12325 => "0000000000000000",12326 => "0000000000000000",
12327 => "0000000000000000",12328 => "0000000000000000",
12329 => "0000000000000000",12330 => "0000000000000000",
12331 => "0000000000000000",12332 => "0000000000000000",
12333 => "0000000000000000",12334 => "0000000000000000",
12335 => "0000000000000000",12336 => "0000000000000000",
12337 => "0000000000000000",12338 => "0000000000000000",
12339 => "0000000000000000",12340 => "0000000000000000",
12341 => "0000000000000000",12342 => "0000000000000000",
12343 => "0000000000000000",12344 => "0000000000000000",
12345 => "0000000000000000",12346 => "0000000000000000",
12347 => "0000000000000000",12348 => "0000000000000000",
12349 => "0000000000000000",12350 => "0000000000000000",
12351 => "0000000000000000",12352 => "0000000000000000",
12353 => "0000000000000000",12354 => "0000000000000000",
12355 => "0000000000000000",12356 => "0000000000000000",
12357 => "0000000000000000",12358 => "0000000000000000",
12359 => "0000000000000000",12360 => "0000000000000000",
12361 => "0000000000000000",12362 => "0000000000000000",
12363 => "0000000000000000",12364 => "0000000000000000",
12365 => "0000000000000000",12366 => "0000000000000000",
12367 => "0000000000000000",12368 => "0000000000000000",
12369 => "0000000000000000",12370 => "0000000000000000",
12371 => "0000000000000000",12372 => "0000000000000000",
12373 => "0000000000000000",12374 => "0000000000000000",
12375 => "0000000000000000",12376 => "0000000000000000",
12377 => "0000000000000000",12378 => "0000000000000000",
12379 => "0000000000000000",12380 => "0000000000000000",
12381 => "0000000000000000",12382 => "0000000000000000",
12383 => "0000000000000000",12384 => "0000000000000000",
12385 => "0000000000000000",12386 => "0000000000000000",
12387 => "0000000000000000",12388 => "0000000000000000",
12389 => "0000000000000000",12390 => "0000000000000000",
12391 => "0000000000000000",12392 => "0000000000000000",
12393 => "0000000000000000",12394 => "0000000000000000",
12395 => "0000000000000000",12396 => "0000000000000000",
12397 => "0000000000000000",12398 => "0000000000000000",
12399 => "0000000000000000",12400 => "0000000000000000",
12401 => "0000000000000000",12402 => "0000000000000000",
12403 => "0000000000000000",12404 => "0000000000000000",
12405 => "0000000000000000",12406 => "0000000000000000",
12407 => "0000000000000000",12408 => "0000000000000000",
12409 => "0000000000000000",12410 => "0000000000000000",
12411 => "0000000000000000",12412 => "0000000000000000",
12413 => "0000000000000000",12414 => "0000000000000000",
12415 => "0000000000000000",12416 => "0000000000000000",
12417 => "0000000000000000",12418 => "0000000000000000",
12419 => "0000000000000000",12420 => "0000000000000000",
12421 => "0000000000000000",12422 => "0000000000000000",
12423 => "0000000000000000",12424 => "0000000000000000",
12425 => "0000000000000000",12426 => "0000000000000000",
12427 => "0000000000000000",12428 => "0000000000000000",
12429 => "0000000000000000",12430 => "0000000000000000",
12431 => "0000000000000000",12432 => "0000000000000000",
12433 => "0000000000000000",12434 => "0000000000000000",
12435 => "0000000000000000",12436 => "0000000000000000",
12437 => "0000000000000000",12438 => "0000000000000000",
12439 => "0000000000000000",12440 => "0000000000000000",
12441 => "0000000000000000",12442 => "0000000000000000",
12443 => "0000000000000000",12444 => "0000000000000000",
12445 => "0000000000000000",12446 => "0000000000000000",
12447 => "0000000000000000",12448 => "0000000000000000",
12449 => "0000000000000000",12450 => "0000000000000000",
12451 => "0000000000000000",12452 => "0000000000000000",
12453 => "0000000000000000",12454 => "0000000000000000",
12455 => "0000000000000000",12456 => "0000000000000000",
12457 => "0000000000000000",12458 => "0000000000000000",
12459 => "0000000000000000",12460 => "0000000000000000",
12461 => "0000000000000000",12462 => "0000000000000000",
12463 => "0000000000000000",12464 => "0000000000000000",
12465 => "0000000000000000",12466 => "0000000000000000",
12467 => "0000000000000000",12468 => "0000000000000000",
12469 => "0000000000000000",12470 => "0000000000000000",
12471 => "0000000000000000",12472 => "0000000000000000",
12473 => "0000000000000000",12474 => "0000000000000000",
12475 => "0000000000000000",12476 => "0000000000000000",
12477 => "0000000000000000",12478 => "0000000000000000",
12479 => "0000000000000000",12480 => "0000000000000000",
12481 => "0000000000000000",12482 => "0000000000000000",
12483 => "0000000000000000",12484 => "0000000000000000",
12485 => "0000000000000000",12486 => "0000000000000000",
12487 => "0000000000000000",12488 => "0000000000000000",
12489 => "0000000000000000",12490 => "0000000000000000",
12491 => "0000000000000000",12492 => "0000000000000000",
12493 => "0000000000000000",12494 => "0000000000000000",
12495 => "0000000000000000",12496 => "0000000000000000",
12497 => "0000000000000000",12498 => "0000000000000000",
12499 => "0000000000000000",12500 => "0000000000000000",
12501 => "0000000000000000",12502 => "0000000000000000",
12503 => "0000000000000000",12504 => "0000000000000000",
12505 => "0000000000000000",12506 => "0000000000000000",
12507 => "0000000000000000",12508 => "0000000000000000",
12509 => "0000000000000000",12510 => "0000000000000000",
12511 => "0000000000000000",12512 => "0000000000000000",
12513 => "0000000000000000",12514 => "0000000000000000",
12515 => "0000000000000000",12516 => "0000000000000000",
12517 => "0000000000000000",12518 => "0000000000000000",
12519 => "0000000000000000",12520 => "0000000000000000",
12521 => "0000000000000000",12522 => "0000000000000000",
12523 => "0000000000000000",12524 => "0000000000000000",
12525 => "0000000000000000",12526 => "0000000000000000",
12527 => "0000000000000000",12528 => "0000000000000000",
12529 => "0000000000000000",12530 => "0000000000000000",
12531 => "0000000000000000",12532 => "0000000000000000",
12533 => "0000000000000000",12534 => "0000000000000000",
12535 => "0000000000000000",12536 => "0000000000000000",
12537 => "0000000000000000",12538 => "0000000000000000",
12539 => "0000000000000000",12540 => "0000000000000000",
12541 => "0000000000000000",12542 => "0000000000000000",
12543 => "0000000000000000",12544 => "0000000000000000",
12545 => "0000000000000000",12546 => "0000000000000000",
12547 => "0000000000000000",12548 => "0000000000000000",
12549 => "0000000000000000",12550 => "0000000000000000",
12551 => "0000000000000000",12552 => "0000000000000000",
12553 => "0000000000000000",12554 => "0000000000000000",
12555 => "0000000000000000",12556 => "0000000000000000",
12557 => "0000000000000000",12558 => "0000000000000000",
12559 => "0000000000000000",12560 => "0000000000000000",
12561 => "0000000000000000",12562 => "0000000000000000",
12563 => "0000000000000000",12564 => "0000000000000000",
12565 => "0000000000000000",12566 => "0000000000000000",
12567 => "0000000000000000",12568 => "0000000000000000",
12569 => "0000000000000000",12570 => "0000000000000000",
12571 => "0000000000000000",12572 => "0000000000000000",
12573 => "0000000000000000",12574 => "0000000000000000",
12575 => "0000000000000000",12576 => "0000000000000000",
12577 => "0000000000000000",12578 => "0000000000000000",
12579 => "0000000000000000",12580 => "0000000000000000",
12581 => "0000000000000000",12582 => "0000000000000000",
12583 => "0000000000000000",12584 => "0000000000000000",
12585 => "0000000000000000",12586 => "0000000000000000",
12587 => "0000000000000000",12588 => "0000000000000000",
12589 => "0000000000000000",12590 => "0000000000000000",
12591 => "0000000000000000",12592 => "0000000000000000",
12593 => "0000000000000000",12594 => "0000000000000000",
12595 => "0000000000000000",12596 => "0000000000000000",
12597 => "0000000000000000",12598 => "0000000000000000",
12599 => "0000000000000000",12600 => "0000000000000000",
12601 => "0000000000000000",12602 => "0000000000000000",
12603 => "0000000000000000",12604 => "0000000000000000",
12605 => "0000000000000000",12606 => "0000000000000000",
12607 => "0000000000000000",12608 => "0000000000000000",
12609 => "0000000000000000",12610 => "0000000000000000",
12611 => "0000000000000000",12612 => "0000000000000000",
12613 => "0000000000000000",12614 => "0000000000000000",
12615 => "0000000000000000",12616 => "0000000000000000",
12617 => "0000000000000000",12618 => "0000000000000000",
12619 => "0000000000000000",12620 => "0000000000000000",
12621 => "0000000000000000",12622 => "0000000000000000",
12623 => "0000000000000000",12624 => "0000000000000000",
12625 => "0000000000000000",12626 => "0000000000000000",
12627 => "0000000000000000",12628 => "0000000000000000",
12629 => "0000000000000000",12630 => "0000000000000000",
12631 => "0000000000000000",12632 => "0000000000000000",
12633 => "0000000000000000",12634 => "0000000000000000",
12635 => "0000000000000000",12636 => "0000000000000000",
12637 => "0000000000000000",12638 => "0000000000000000",
12639 => "0000000000000000",12640 => "0000000000000000",
12641 => "0000000000000000",12642 => "0000000000000000",
12643 => "0000000000000000",12644 => "0000000000000000",
12645 => "0000000000000000",12646 => "0000000000000000",
12647 => "0000000000000000",12648 => "0000000000000000",
12649 => "0000000000000000",12650 => "0000000000000000",
12651 => "0000000000000000",12652 => "0000000000000000",
12653 => "0000000000000000",12654 => "0000000000000000",
12655 => "0000000000000000",12656 => "0000000000000000",
12657 => "0000000000000000",12658 => "0000000000000000",
12659 => "0000000000000000",12660 => "0000000000000000",
12661 => "0000000000000000",12662 => "0000000000000000",
12663 => "0000000000000000",12664 => "0000000000000000",
12665 => "0000000000000000",12666 => "0000000000000000",
12667 => "0000000000000000",12668 => "0000000000000000",
12669 => "0000000000000000",12670 => "0000000000000000",
12671 => "0000000000000000",12672 => "0000000000000000",
12673 => "0000000000000000",12674 => "0000000000000000",
12675 => "0000000000000000",12676 => "0000000000000000",
12677 => "0000000000000000",12678 => "0000000000000000",
12679 => "0000000000000000",12680 => "0000000000000000",
12681 => "0000000000000000",12682 => "0000000000000000",
12683 => "0000000000000000",12684 => "0000000000000000",
12685 => "0000000000000000",12686 => "0000000000000000",
12687 => "0000000000000000",12688 => "0000000000000000",
12689 => "0000000000000000",12690 => "0000000000000000",
12691 => "0000000000000000",12692 => "0000000000000000",
12693 => "0000000000000000",12694 => "0000000000000000",
12695 => "0000000000000000",12696 => "0000000000000000",
12697 => "0000000000000000",12698 => "0000000000000000",
12699 => "0000000000000000",12700 => "0000000000000000",
12701 => "0000000000000000",12702 => "0000000000000000",
12703 => "0000000000000000",12704 => "0000000000000000",
12705 => "0000000000000000",12706 => "0000000000000000",
12707 => "0000000000000000",12708 => "0000000000000000",
12709 => "0000000000000000",12710 => "0000000000000000",
12711 => "0000000000000000",12712 => "0000000000000000",
12713 => "0000000000000000",12714 => "0000000000000000",
12715 => "0000000000000000",12716 => "0000000000000000",
12717 => "0000000000000000",12718 => "0000000000000000",
12719 => "0000000000000000",12720 => "0000000000000000",
12721 => "0000000000000000",12722 => "0000000000000000",
12723 => "0000000000000000",12724 => "0000000000000000",
12725 => "0000000000000000",12726 => "0000000000000000",
12727 => "0000000000000000",12728 => "0000000000000000",
12729 => "0000000000000000",12730 => "0000000000000000",
12731 => "0000000000000000",12732 => "0000000000000000",
12733 => "0000000000000000",12734 => "0000000000000000",
12735 => "0000000000000000",12736 => "0000000000000000",
12737 => "0000000000000000",12738 => "0000000000000000",
12739 => "0000000000000000",12740 => "0000000000000000",
12741 => "0000000000000000",12742 => "0000000000000000",
12743 => "0000000000000000",12744 => "0000000000000000",
12745 => "0000000000000000",12746 => "0000000000000000",
12747 => "0000000000000000",12748 => "0000000000000000",
12749 => "0000000000000000",12750 => "0000000000000000",
12751 => "0000000000000000",12752 => "0000000000000000",
12753 => "0000000000000000",12754 => "0000000000000000",
12755 => "0000000000000000",12756 => "0000000000000000",
12757 => "0000000000000000",12758 => "0000000000000000",
12759 => "0000000000000000",12760 => "0000000000000000",
12761 => "0000000000000000",12762 => "0000000000000000",
12763 => "0000000000000000",12764 => "0000000000000000",
12765 => "0000000000000000",12766 => "0000000000000000",
12767 => "0000000000000000",12768 => "0000000000000000",
12769 => "0000000000000000",12770 => "0000000000000000",
12771 => "0000000000000000",12772 => "0000000000000000",
12773 => "0000000000000000",12774 => "0000000000000000",
12775 => "0000000000000000",12776 => "0000000000000000",
12777 => "0000000000000000",12778 => "0000000000000000",
12779 => "0000000000000000",12780 => "0000000000000000",
12781 => "0000000000000000",12782 => "0000000000000000",
12783 => "0000000000000000",12784 => "0000000000000000",
12785 => "0000000000000000",12786 => "0000000000000000",
12787 => "0000000000000000",12788 => "0000000000000000",
12789 => "0000000000000000",12790 => "0000000000000000",
12791 => "0000000000000000",12792 => "0000000000000000",
12793 => "0000000000000000",12794 => "0000000000000000",
12795 => "0000000000000000",12796 => "0000000000000000",
12797 => "0000000000000000",12798 => "0000000000000000",
12799 => "0000000000000000",12800 => "0000000000000000",
12801 => "0000000000000000",12802 => "0000000000000000",
12803 => "0000000000000000",12804 => "0000000000000000",
12805 => "0000000000000000",12806 => "0000000000000000",
12807 => "0000000000000000",12808 => "0000000000000000",
12809 => "0000000000000000",12810 => "0000000000000000",
12811 => "0000000000000000",12812 => "0000000000000000",
12813 => "0000000000000000",12814 => "0000000000000000",
12815 => "0000000000000000",12816 => "0000000000000000",
12817 => "0000000000000000",12818 => "0000000000000000",
12819 => "0000000000000000",12820 => "0000000000000000",
12821 => "0000000000000000",12822 => "0000000000000000",
12823 => "0000000000000000",12824 => "0000000000000000",
12825 => "0000000000000000",12826 => "0000000000000000",
12827 => "0000000000000000",12828 => "0000000000000000",
12829 => "0000000000000000",12830 => "0000000000000000",
12831 => "0000000000000000",12832 => "0000000000000000",
12833 => "0000000000000000",12834 => "0000000000000000",
12835 => "0000000000000000",12836 => "0000000000000000",
12837 => "0000000000000000",12838 => "0000000000000000",
12839 => "0000000000000000",12840 => "0000000000000000",
12841 => "0000000000000000",12842 => "0000000000000000",
12843 => "0000000000000000",12844 => "0000000000000000",
12845 => "0000000000000000",12846 => "0000000000000000",
12847 => "0000000000000000",12848 => "0000000000000000",
12849 => "0000000000000000",12850 => "0000000000000000",
12851 => "0000000000000000",12852 => "0000000000000000",
12853 => "0000000000000000",12854 => "0000000000000000",
12855 => "0000000000000000",12856 => "0000000000000000",
12857 => "0000000000000000",12858 => "0000000000000000",
12859 => "0000000000000000",12860 => "0000000000000000",
12861 => "0000000000000000",12862 => "0000000000000000",
12863 => "0000000000000000",12864 => "0000000000000000",
12865 => "0000000000000000",12866 => "0000000000000000",
12867 => "0000000000000000",12868 => "0000000000000000",
12869 => "0000000000000000",12870 => "0000000000000000",
12871 => "0000000000000000",12872 => "0000000000000000",
12873 => "0000000000000000",12874 => "0000000000000000",
12875 => "0000000000000000",12876 => "0000000000000000",
12877 => "0000000000000000",12878 => "0000000000000000",
12879 => "0000000000000000",12880 => "0000000000000000",
12881 => "0000000000000000",12882 => "0000000000000000",
12883 => "0000000000000000",12884 => "0000000000000000",
12885 => "0000000000000000",12886 => "0000000000000000",
12887 => "0000000000000000",12888 => "0000000000000000",
12889 => "0000000000000000",12890 => "0000000000000000",
12891 => "0000000000000000",12892 => "0000000000000000",
12893 => "0000000000000000",12894 => "0000000000000000",
12895 => "0000000000000000",12896 => "0000000000000000",
12897 => "0000000000000000",12898 => "0000000000000000",
12899 => "0000000000000000",12900 => "0000000000000000",
12901 => "0000000000000000",12902 => "0000000000000000",
12903 => "0000000000000000",12904 => "0000000000000000",
12905 => "0000000000000000",12906 => "0000000000000000",
12907 => "0000000000000000",12908 => "0000000000000000",
12909 => "0000000000000000",12910 => "0000000000000000",
12911 => "0000000000000000",12912 => "0000000000000000",
12913 => "0000000000000000",12914 => "0000000000000000",
12915 => "0000000000000000",12916 => "0000000000000000",
12917 => "0000000000000000",12918 => "0000000000000000",
12919 => "0000000000000000",12920 => "0000000000000000",
12921 => "0000000000000000",12922 => "0000000000000000",
12923 => "0000000000000000",12924 => "0000000000000000",
12925 => "0000000000000000",12926 => "0000000000000000",
12927 => "0000000000000000",12928 => "0000000000000000",
12929 => "0000000000000000",12930 => "0000000000000000",
12931 => "0000000000000000",12932 => "0000000000000000",
12933 => "0000000000000000",12934 => "0000000000000000",
12935 => "0000000000000000",12936 => "0000000000000000",
12937 => "0000000000000000",12938 => "0000000000000000",
12939 => "0000000000000000",12940 => "0000000000000000",
12941 => "0000000000000000",12942 => "0000000000000000",
12943 => "0000000000000000",12944 => "0000000000000000",
12945 => "0000000000000000",12946 => "0000000000000000",
12947 => "0000000000000000",12948 => "0000000000000000",
12949 => "0000000000000000",12950 => "0000000000000000",
12951 => "0000000000000000",12952 => "0000000000000000",
12953 => "0000000000000000",12954 => "0000000000000000",
12955 => "0000000000000000",12956 => "0000000000000000",
12957 => "0000000000000000",12958 => "0000000000000000",
12959 => "0000000000000000",12960 => "0000000000000000",
12961 => "0000000000000000",12962 => "0000000000000000",
12963 => "0000000000000000",12964 => "0000000000000000",
12965 => "0000000000000000",12966 => "0000000000000000",
12967 => "0000000000000000",12968 => "0000000000000000",
12969 => "0000000000000000",12970 => "0000000000000000",
12971 => "0000000000000000",12972 => "0000000000000000",
12973 => "0000000000000000",12974 => "0000000000000000",
12975 => "0000000000000000",12976 => "0000000000000000",
12977 => "0000000000000000",12978 => "0000000000000000",
12979 => "0000000000000000",12980 => "0000000000000000",
12981 => "0000000000000000",12982 => "0000000000000000",
12983 => "0000000000000000",12984 => "0000000000000000",
12985 => "0000000000000000",12986 => "0000000000000000",
12987 => "0000000000000000",12988 => "0000000000000000",
12989 => "0000000000000000",12990 => "0000000000000000",
12991 => "0000000000000000",12992 => "0000000000000000",
12993 => "0000000000000000",12994 => "0000000000000000",
12995 => "0000000000000000",12996 => "0000000000000000",
12997 => "0000000000000000",12998 => "0000000000000000",
12999 => "0000000000000000",13000 => "0000000000000000",
13001 => "0000000000000000",13002 => "0000000000000000",
13003 => "0000000000000000",13004 => "0000000000000000",
13005 => "0000000000000000",13006 => "0000000000000000",
13007 => "0000000000000000",13008 => "0000000000000000",
13009 => "0000000000000000",13010 => "0000000000000000",
13011 => "0000000000000000",13012 => "0000000000000000",
13013 => "0000000000000000",13014 => "0000000000000000",
13015 => "0000000000000000",13016 => "0000000000000000",
13017 => "0000000000000000",13018 => "0000000000000000",
13019 => "0000000000000000",13020 => "0000000000000000",
13021 => "0000000000000000",13022 => "0000000000000000",
13023 => "0000000000000000",13024 => "0000000000000000",
13025 => "0000000000000000",13026 => "0000000000000000",
13027 => "0000000000000000",13028 => "0000000000000000",
13029 => "0000000000000000",13030 => "0000000000000000",
13031 => "0000000000000000",13032 => "0000000000000000",
13033 => "0000000000000000",13034 => "0000000000000000",
13035 => "0000000000000000",13036 => "0000000000000000",
13037 => "0000000000000000",13038 => "0000000000000000",
13039 => "0000000000000000",13040 => "0000000000000000",
13041 => "0000000000000000",13042 => "0000000000000000",
13043 => "0000000000000000",13044 => "0000000000000000",
13045 => "0000000000000000",13046 => "0000000000000000",
13047 => "0000000000000000",13048 => "0000000000000000",
13049 => "0000000000000000",13050 => "0000000000000000",
13051 => "0000000000000000",13052 => "0000000000000000",
13053 => "0000000000000000",13054 => "0000000000000000",
13055 => "0000000000000000",13056 => "0000000000000000",
13057 => "0000000000000000",13058 => "0000000000000000",
13059 => "0000000000000000",13060 => "0000000000000000",
13061 => "0000000000000000",13062 => "0000000000000000",
13063 => "0000000000000000",13064 => "0000000000000000",
13065 => "0000000000000000",13066 => "0000000000000000",
13067 => "0000000000000000",13068 => "0000000000000000",
13069 => "0000000000000000",13070 => "0000000000000000",
13071 => "0000000000000000",13072 => "0000000000000000",
13073 => "0000000000000000",13074 => "0000000000000000",
13075 => "0000000000000000",13076 => "0000000000000000",
13077 => "0000000000000000",13078 => "0000000000000000",
13079 => "0000000000000000",13080 => "0000000000000000",
13081 => "0000000000000000",13082 => "0000000000000000",
13083 => "0000000000000000",13084 => "0000000000000000",
13085 => "0000000000000000",13086 => "0000000000000000",
13087 => "0000000000000000",13088 => "0000000000000000",
13089 => "0000000000000000",13090 => "0000000000000000",
13091 => "0000000000000000",13092 => "0000000000000000",
13093 => "0000000000000000",13094 => "0000000000000000",
13095 => "0000000000000000",13096 => "0000000000000000",
13097 => "0000000000000000",13098 => "0000000000000000",
13099 => "0000000000000000",13100 => "0000000000000000",
13101 => "0000000000000000",13102 => "0000000000000000",
13103 => "0000000000000000",13104 => "0000000000000000",
13105 => "0000000000000000",13106 => "0000000000000000",
13107 => "0000000000000000",13108 => "0000000000000000",
13109 => "0000000000000000",13110 => "0000000000000000",
13111 => "0000000000000000",13112 => "0000000000000000",
13113 => "0000000000000000",13114 => "0000000000000000",
13115 => "0000000000000000",13116 => "0000000000000000",
13117 => "0000000000000000",13118 => "0000000000000000",
13119 => "0000000000000000",13120 => "0000000000000000",
13121 => "0000000000000000",13122 => "0000000000000000",
13123 => "0000000000000000",13124 => "0000000000000000",
13125 => "0000000000000000",13126 => "0000000000000000",
13127 => "0000000000000000",13128 => "0000000000000000",
13129 => "0000000000000000",13130 => "0000000000000000",
13131 => "0000000000000000",13132 => "0000000000000000",
13133 => "0000000000000000",13134 => "0000000000000000",
13135 => "0000000000000000",13136 => "0000000000000000",
13137 => "0000000000000000",13138 => "0000000000000000",
13139 => "0000000000000000",13140 => "0000000000000000",
13141 => "0000000000000000",13142 => "0000000000000000",
13143 => "0000000000000000",13144 => "0000000000000000",
13145 => "0000000000000000",13146 => "0000000000000000",
13147 => "0000000000000000",13148 => "0000000000000000",
13149 => "0000000000000000",13150 => "0000000000000000",
13151 => "0000000000000000",13152 => "0000000000000000",
13153 => "0000000000000000",13154 => "0000000000000000",
13155 => "0000000000000000",13156 => "0000000000000000",
13157 => "0000000000000000",13158 => "0000000000000000",
13159 => "0000000000000000",13160 => "0000000000000000",
13161 => "0000000000000000",13162 => "0000000000000000",
13163 => "0000000000000000",13164 => "0000000000000000",
13165 => "0000000000000000",13166 => "0000000000000000",
13167 => "0000000000000000",13168 => "0000000000000000",
13169 => "0000000000000000",13170 => "0000000000000000",
13171 => "0000000000000000",13172 => "0000000000000000",
13173 => "0000000000000000",13174 => "0000000000000000",
13175 => "0000000000000000",13176 => "0000000000000000",
13177 => "0000000000000000",13178 => "0000000000000000",
13179 => "0000000000000000",13180 => "0000000000000000",
13181 => "0000000000000000",13182 => "0000000000000000",
13183 => "0000000000000000",13184 => "0000000000000000",
13185 => "0000000000000000",13186 => "0000000000000000",
13187 => "0000000000000000",13188 => "0000000000000000",
13189 => "0000000000000000",13190 => "0000000000000000",
13191 => "0000000000000000",13192 => "0000000000000000",
13193 => "0000000000000000",13194 => "0000000000000000",
13195 => "0000000000000000",13196 => "0000000000000000",
13197 => "0000000000000000",13198 => "0000000000000000",
13199 => "0000000000000000",13200 => "0000000000000000",
13201 => "0000000000000000",13202 => "0000000000000000",
13203 => "0000000000000000",13204 => "0000000000000000",
13205 => "0000000000000000",13206 => "0000000000000000",
13207 => "0000000000000000",13208 => "0000000000000000",
13209 => "0000000000000000",13210 => "0000000000000000",
13211 => "0000000000000000",13212 => "0000000000000000",
13213 => "0000000000000000",13214 => "0000000000000000",
13215 => "0000000000000000",13216 => "0000000000000000",
13217 => "0000000000000000",13218 => "0000000000000000",
13219 => "0000000000000000",13220 => "0000000000000000",
13221 => "0000000000000000",13222 => "0000000000000000",
13223 => "0000000000000000",13224 => "0000000000000000",
13225 => "0000000000000000",13226 => "0000000000000000",
13227 => "0000000000000000",13228 => "0000000000000000",
13229 => "0000000000000000",13230 => "0000000000000000",
13231 => "0000000000000000",13232 => "0000000000000000",
13233 => "0000000000000000",13234 => "0000000000000000",
13235 => "0000000000000000",13236 => "0000000000000000",
13237 => "0000000000000000",13238 => "0000000000000000",
13239 => "0000000000000000",13240 => "0000000000000000",
13241 => "0000000000000000",13242 => "0000000000000000",
13243 => "0000000000000000",13244 => "0000000000000000",
13245 => "0000000000000000",13246 => "0000000000000000",
13247 => "0000000000000000",13248 => "0000000000000000",
13249 => "0000000000000000",13250 => "0000000000000000",
13251 => "0000000000000000",13252 => "0000000000000000",
13253 => "0000000000000000",13254 => "0000000000000000",
13255 => "0000000000000000",13256 => "0000000000000000",
13257 => "0000000000000000",13258 => "0000000000000000",
13259 => "0000000000000000",13260 => "0000000000000000",
13261 => "0000000000000000",13262 => "0000000000000000",
13263 => "0000000000000000",13264 => "0000000000000000",
13265 => "0000000000000000",13266 => "0000000000000000",
13267 => "0000000000000000",13268 => "0000000000000000",
13269 => "0000000000000000",13270 => "0000000000000000",
13271 => "0000000000000000",13272 => "0000000000000000",
13273 => "0000000000000000",13274 => "0000000000000000",
13275 => "0000000000000000",13276 => "0000000000000000",
13277 => "0000000000000000",13278 => "0000000000000000",
13279 => "0000000000000000",13280 => "0000000000000000",
13281 => "0000000000000000",13282 => "0000000000000000",
13283 => "0000000000000000",13284 => "0000000000000000",
13285 => "0000000000000000",13286 => "0000000000000000",
13287 => "0000000000000000",13288 => "0000000000000000",
13289 => "0000000000000000",13290 => "0000000000000000",
13291 => "0000000000000000",13292 => "0000000000000000",
13293 => "0000000000000000",13294 => "0000000000000000",
13295 => "0000000000000000",13296 => "0000000000000000",
13297 => "0000000000000000",13298 => "0000000000000000",
13299 => "0000000000000000",13300 => "0000000000000000",
13301 => "0000000000000000",13302 => "0000000000000000",
13303 => "0000000000000000",13304 => "0000000000000000",
13305 => "0000000000000000",13306 => "0000000000000000",
13307 => "0000000000000000",13308 => "0000000000000000",
13309 => "0000000000000000",13310 => "0000000000000000",
13311 => "0000000000000000",13312 => "0000000000000000",
13313 => "0000000000000000",13314 => "0000000000000000",
13315 => "0000000000000000",13316 => "0000000000000000",
13317 => "0000000000000000",13318 => "0000000000000000",
13319 => "0000000000000000",13320 => "0000000000000000",
13321 => "0000000000000000",13322 => "0000000000000000",
13323 => "0000000000000000",13324 => "0000000000000000",
13325 => "0000000000000000",13326 => "0000000000000000",
13327 => "0000000000000000",13328 => "0000000000000000",
13329 => "0000000000000000",13330 => "0000000000000000",
13331 => "0000000000000000",13332 => "0000000000000000",
13333 => "0000000000000000",13334 => "0000000000000000",
13335 => "0000000000000000",13336 => "0000000000000000",
13337 => "0000000000000000",13338 => "0000000000000000",
13339 => "0000000000000000",13340 => "0000000000000000",
13341 => "0000000000000000",13342 => "0000000000000000",
13343 => "0000000000000000",13344 => "0000000000000000",
13345 => "0000000000000000",13346 => "0000000000000000",
13347 => "0000000000000000",13348 => "0000000000000000",
13349 => "0000000000000000",13350 => "0000000000000000",
13351 => "0000000000000000",13352 => "0000000000000000",
13353 => "0000000000000000",13354 => "0000000000000000",
13355 => "0000000000000000",13356 => "0000000000000000",
13357 => "0000000000000000",13358 => "0000000000000000",
13359 => "0000000000000000",13360 => "0000000000000000",
13361 => "0000000000000000",13362 => "0000000000000000",
13363 => "0000000000000000",13364 => "0000000000000000",
13365 => "0000000000000000",13366 => "0000000000000000",
13367 => "0000000000000000",13368 => "0000000000000000",
13369 => "0000000000000000",13370 => "0000000000000000",
13371 => "0000000000000000",13372 => "0000000000000000",
13373 => "0000000000000000",13374 => "0000000000000000",
13375 => "0000000000000000",13376 => "0000000000000000",
13377 => "0000000000000000",13378 => "0000000000000000",
13379 => "0000000000000000",13380 => "0000000000000000",
13381 => "0000000000000000",13382 => "0000000000000000",
13383 => "0000000000000000",13384 => "0000000000000000",
13385 => "0000000000000000",13386 => "0000000000000000",
13387 => "0000000000000000",13388 => "0000000000000000",
13389 => "0000000000000000",13390 => "0000000000000000",
13391 => "0000000000000000",13392 => "0000000000000000",
13393 => "0000000000000000",13394 => "0000000000000000",
13395 => "0000000000000000",13396 => "0000000000000000",
13397 => "0000000000000000",13398 => "0000000000000000",
13399 => "0000000000000000",13400 => "0000000000000000",
13401 => "0000000000000000",13402 => "0000000000000000",
13403 => "0000000000000000",13404 => "0000000000000000",
13405 => "0000000000000000",13406 => "0000000000000000",
13407 => "0000000000000000",13408 => "0000000000000000",
13409 => "0000000000000000",13410 => "0000000000000000",
13411 => "0000000000000000",13412 => "0000000000000000",
13413 => "0000000000000000",13414 => "0000000000000000",
13415 => "0000000000000000",13416 => "0000000000000000",
13417 => "0000000000000000",13418 => "0000000000000000",
13419 => "0000000000000000",13420 => "0000000000000000",
13421 => "0000000000000000",13422 => "0000000000000000",
13423 => "0000000000000000",13424 => "0000000000000000",
13425 => "0000000000000000",13426 => "0000000000000000",
13427 => "0000000000000000",13428 => "0000000000000000",
13429 => "0000000000000000",13430 => "0000000000000000",
13431 => "0000000000000000",13432 => "0000000000000000",
13433 => "0000000000000000",13434 => "0000000000000000",
13435 => "0000000000000000",13436 => "0000000000000000",
13437 => "0000000000000000",13438 => "0000000000000000",
13439 => "0000000000000000",13440 => "0000000000000000",
13441 => "0000000000000000",13442 => "0000000000000000",
13443 => "0000000000000000",13444 => "0000000000000000",
13445 => "0000000000000000",13446 => "0000000000000000",
13447 => "0000000000000000",13448 => "0000000000000000",
13449 => "0000000000000000",13450 => "0000000000000000",
13451 => "0000000000000000",13452 => "0000000000000000",
13453 => "0000000000000000",13454 => "0000000000000000",
13455 => "0000000000000000",13456 => "0000000000000000",
13457 => "0000000000000000",13458 => "0000000000000000",
13459 => "0000000000000000",13460 => "0000000000000000",
13461 => "0000000000000000",13462 => "0000000000000000",
13463 => "0000000000000000",13464 => "0000000000000000",
13465 => "0000000000000000",13466 => "0000000000000000",
13467 => "0000000000000000",13468 => "0000000000000000",
13469 => "0000000000000000",13470 => "0000000000000000",
13471 => "0000000000000000",13472 => "0000000000000000",
13473 => "0000000000000000",13474 => "0000000000000000",
13475 => "0000000000000000",13476 => "0000000000000000",
13477 => "0000000000000000",13478 => "0000000000000000",
13479 => "0000000000000000",13480 => "0000000000000000",
13481 => "0000000000000000",13482 => "0000000000000000",
13483 => "0000000000000000",13484 => "0000000000000000",
13485 => "0000000000000000",13486 => "0000000000000000",
13487 => "0000000000000000",13488 => "0000000000000000",
13489 => "0000000000000000",13490 => "0000000000000000",
13491 => "0000000000000000",13492 => "0000000000000000",
13493 => "0000000000000000",13494 => "0000000000000000",
13495 => "0000000000000000",13496 => "0000000000000000",
13497 => "0000000000000000",13498 => "0000000000000000",
13499 => "0000000000000000",13500 => "0000000000000000",
13501 => "0000000000000000",13502 => "0000000000000000",
13503 => "0000000000000000",13504 => "0000000000000000",
13505 => "0000000000000000",13506 => "0000000000000000",
13507 => "0000000000000000",13508 => "0000000000000000",
13509 => "0000000000000000",13510 => "0000000000000000",
13511 => "0000000000000000",13512 => "0000000000000000",
13513 => "0000000000000000",13514 => "0000000000000000",
13515 => "0000000000000000",13516 => "0000000000000000",
13517 => "0000000000000000",13518 => "0000000000000000",
13519 => "0000000000000000",13520 => "0000000000000000",
13521 => "0000000000000000",13522 => "0000000000000000",
13523 => "0000000000000000",13524 => "0000000000000000",
13525 => "0000000000000000",13526 => "0000000000000000",
13527 => "0000000000000000",13528 => "0000000000000000",
13529 => "0000000000000000",13530 => "0000000000000000",
13531 => "0000000000000000",13532 => "0000000000000000",
13533 => "0000000000000000",13534 => "0000000000000000",
13535 => "0000000000000000",13536 => "0000000000000000",
13537 => "0000000000000000",13538 => "0000000000000000",
13539 => "0000000000000000",13540 => "0000000000000000",
13541 => "0000000000000000",13542 => "0000000000000000",
13543 => "0000000000000000",13544 => "0000000000000000",
13545 => "0000000000000000",13546 => "0000000000000000",
13547 => "0000000000000000",13548 => "0000000000000000",
13549 => "0000000000000000",13550 => "0000000000000000",
13551 => "0000000000000000",13552 => "0000000000000000",
13553 => "0000000000000000",13554 => "0000000000000000",
13555 => "0000000000000000",13556 => "0000000000000000",
13557 => "0000000000000000",13558 => "0000000000000000",
13559 => "0000000000000000",13560 => "0000000000000000",
13561 => "0000000000000000",13562 => "0000000000000000",
13563 => "0000000000000000",13564 => "0000000000000000",
13565 => "0000000000000000",13566 => "0000000000000000",
13567 => "0000000000000000",13568 => "0000000000000000",
13569 => "0000000000000000",13570 => "0000000000000000",
13571 => "0000000000000000",13572 => "0000000000000000",
13573 => "0000000000000000",13574 => "0000000000000000",
13575 => "0000000000000000",13576 => "0000000000000000",
13577 => "0000000000000000",13578 => "0000000000000000",
13579 => "0000000000000000",13580 => "0000000000000000",
13581 => "0000000000000000",13582 => "0000000000000000",
13583 => "0000000000000000",13584 => "0000000000000000",
13585 => "0000000000000000",13586 => "0000000000000000",
13587 => "0000000000000000",13588 => "0000000000000000",
13589 => "0000000000000000",13590 => "0000000000000000",
13591 => "0000000000000000",13592 => "0000000000000000",
13593 => "0000000000000000",13594 => "0000000000000000",
13595 => "0000000000000000",13596 => "0000000000000000",
13597 => "0000000000000000",13598 => "0000000000000000",
13599 => "0000000000000000",13600 => "0000000000000000",
13601 => "0000000000000000",13602 => "0000000000000000",
13603 => "0000000000000000",13604 => "0000000000000000",
13605 => "0000000000000000",13606 => "0000000000000000",
13607 => "0000000000000000",13608 => "0000000000000000",
13609 => "0000000000000000",13610 => "0000000000000000",
13611 => "0000000000000000",13612 => "0000000000000000",
13613 => "0000000000000000",13614 => "0000000000000000",
13615 => "0000000000000000",13616 => "0000000000000000",
13617 => "0000000000000000",13618 => "0000000000000000",
13619 => "0000000000000000",13620 => "0000000000000000",
13621 => "0000000000000000",13622 => "0000000000000000",
13623 => "0000000000000000",13624 => "0000000000000000",
13625 => "0000000000000000",13626 => "0000000000000000",
13627 => "0000000000000000",13628 => "0000000000000000",
13629 => "0000000000000000",13630 => "0000000000000000",
13631 => "0000000000000000",13632 => "0000000000000000",
13633 => "0000000000000000",13634 => "0000000000000000",
13635 => "0000000000000000",13636 => "0000000000000000",
13637 => "0000000000000000",13638 => "0000000000000000",
13639 => "0000000000000000",13640 => "0000000000000000",
13641 => "0000000000000000",13642 => "0000000000000000",
13643 => "0000000000000000",13644 => "0000000000000000",
13645 => "0000000000000000",13646 => "0000000000000000",
13647 => "0000000000000000",13648 => "0000000000000000",
13649 => "0000000000000000",13650 => "0000000000000000",
13651 => "0000000000000000",13652 => "0000000000000000",
13653 => "0000000000000000",13654 => "0000000000000000",
13655 => "0000000000000000",13656 => "0000000000000000",
13657 => "0000000000000000",13658 => "0000000000000000",
13659 => "0000000000000000",13660 => "0000000000000000",
13661 => "0000000000000000",13662 => "0000000000000000",
13663 => "0000000000000000",13664 => "0000000000000000",
13665 => "0000000000000000",13666 => "0000000000000000",
13667 => "0000000000000000",13668 => "0000000000000000",
13669 => "0000000000000000",13670 => "0000000000000000",
13671 => "0000000000000000",13672 => "0000000000000000",
13673 => "0000000000000000",13674 => "0000000000000000",
13675 => "0000000000000000",13676 => "0000000000000000",
13677 => "0000000000000000",13678 => "0000000000000000",
13679 => "0000000000000000",13680 => "0000000000000000",
13681 => "0000000000000000",13682 => "0000000000000000",
13683 => "0000000000000000",13684 => "0000000000000000",
13685 => "0000000000000000",13686 => "0000000000000000",
13687 => "0000000000000000",13688 => "0000000000000000",
13689 => "0000000000000000",13690 => "0000000000000000",
13691 => "0000000000000000",13692 => "0000000000000000",
13693 => "0000000000000000",13694 => "0000000000000000",
13695 => "0000000000000000",13696 => "0000000000000000",
13697 => "0000000000000000",13698 => "0000000000000000",
13699 => "0000000000000000",13700 => "0000000000000000",
13701 => "0000000000000000",13702 => "0000000000000000",
13703 => "0000000000000000",13704 => "0000000000000000",
13705 => "0000000000000000",13706 => "0000000000000000",
13707 => "0000000000000000",13708 => "0000000000000000",
13709 => "0000000000000000",13710 => "0000000000000000",
13711 => "0000000000000000",13712 => "0000000000000000",
13713 => "0000000000000000",13714 => "0000000000000000",
13715 => "0000000000000000",13716 => "0000000000000000",
13717 => "0000000000000000",13718 => "0000000000000000",
13719 => "0000000000000000",13720 => "0000000000000000",
13721 => "0000000000000000",13722 => "0000000000000000",
13723 => "0000000000000000",13724 => "0000000000000000",
13725 => "0000000000000000",13726 => "0000000000000000",
13727 => "0000000000000000",13728 => "0000000000000000",
13729 => "0000000000000000",13730 => "0000000000000000",
13731 => "0000000000000000",13732 => "0000000000000000",
13733 => "0000000000000000",13734 => "0000000000000000",
13735 => "0000000000000000",13736 => "0000000000000000",
13737 => "0000000000000000",13738 => "0000000000000000",
13739 => "0000000000000000",13740 => "0000000000000000",
13741 => "0000000000000000",13742 => "0000000000000000",
13743 => "0000000000000000",13744 => "0000000000000000",
13745 => "0000000000000000",13746 => "0000000000000000",
13747 => "0000000000000000",13748 => "0000000000000000",
13749 => "0000000000000000",13750 => "0000000000000000",
13751 => "0000000000000000",13752 => "0000000000000000",
13753 => "0000000000000000",13754 => "0000000000000000",
13755 => "0000000000000000",13756 => "0000000000000000",
13757 => "0000000000000000",13758 => "0000000000000000",
13759 => "0000000000000000",13760 => "0000000000000000",
13761 => "0000000000000000",13762 => "0000000000000000",
13763 => "0000000000000000",13764 => "0000000000000000",
13765 => "0000000000000000",13766 => "0000000000000000",
13767 => "0000000000000000",13768 => "0000000000000000",
13769 => "0000000000000000",13770 => "0000000000000000",
13771 => "0000000000000000",13772 => "0000000000000000",
13773 => "0000000000000000",13774 => "0000000000000000",
13775 => "0000000000000000",13776 => "0000000000000000",
13777 => "0000000000000000",13778 => "0000000000000000",
13779 => "0000000000000000",13780 => "0000000000000000",
13781 => "0000000000000000",13782 => "0000000000000000",
13783 => "0000000000000000",13784 => "0000000000000000",
13785 => "0000000000000000",13786 => "0000000000000000",
13787 => "0000000000000000",13788 => "0000000000000000",
13789 => "0000000000000000",13790 => "0000000000000000",
13791 => "0000000000000000",13792 => "0000000000000000",
13793 => "0000000000000000",13794 => "0000000000000000",
13795 => "0000000000000000",13796 => "0000000000000000",
13797 => "0000000000000000",13798 => "0000000000000000",
13799 => "0000000000000000",13800 => "0000000000000000",
13801 => "0000000000000000",13802 => "0000000000000000",
13803 => "0000000000000000",13804 => "0000000000000000",
13805 => "0000000000000000",13806 => "0000000000000000",
13807 => "0000000000000000",13808 => "0000000000000000",
13809 => "0000000000000000",13810 => "0000000000000000",
13811 => "0000000000000000",13812 => "0000000000000000",
13813 => "0000000000000000",13814 => "0000000000000000",
13815 => "0000000000000000",13816 => "0000000000000000",
13817 => "0000000000000000",13818 => "0000000000000000",
13819 => "0000000000000000",13820 => "0000000000000000",
13821 => "0000000000000000",13822 => "0000000000000000",
13823 => "0000000000000000",13824 => "0000000000000000",
13825 => "0000000000000000",13826 => "0000000000000000",
13827 => "0000000000000000",13828 => "0000000000000000",
13829 => "0000000000000000",13830 => "0000000000000000",
13831 => "0000000000000000",13832 => "0000000000000000",
13833 => "0000000000000000",13834 => "0000000000000000",
13835 => "0000000000000000",13836 => "0000000000000000",
13837 => "0000000000000000",13838 => "0000000000000000",
13839 => "0000000000000000",13840 => "0000000000000000",
13841 => "0000000000000000",13842 => "0000000000000000",
13843 => "0000000000000000",13844 => "0000000000000000",
13845 => "0000000000000000",13846 => "0000000000000000",
13847 => "0000000000000000",13848 => "0000000000000000",
13849 => "0000000000000000",13850 => "0000000000000000",
13851 => "0000000000000000",13852 => "0000000000000000",
13853 => "0000000000000000",13854 => "0000000000000000",
13855 => "0000000000000000",13856 => "0000000000000000",
13857 => "0000000000000000",13858 => "0000000000000000",
13859 => "0000000000000000",13860 => "0000000000000000",
13861 => "0000000000000000",13862 => "0000000000000000",
13863 => "0000000000000000",13864 => "0000000000000000",
13865 => "0000000000000000",13866 => "0000000000000000",
13867 => "0000000000000000",13868 => "0000000000000000",
13869 => "0000000000000000",13870 => "0000000000000000",
13871 => "0000000000000000",13872 => "0000000000000000",
13873 => "0000000000000000",13874 => "0000000000000000",
13875 => "0000000000000000",13876 => "0000000000000000",
13877 => "0000000000000000",13878 => "0000000000000000",
13879 => "0000000000000000",13880 => "0000000000000000",
13881 => "0000000000000000",13882 => "0000000000000000",
13883 => "0000000000000000",13884 => "0000000000000000",
13885 => "0000000000000000",13886 => "0000000000000000",
13887 => "0000000000000000",13888 => "0000000000000000",
13889 => "0000000000000000",13890 => "0000000000000000",
13891 => "0000000000000000",13892 => "0000000000000000",
13893 => "0000000000000000",13894 => "0000000000000000",
13895 => "0000000000000000",13896 => "0000000000000000",
13897 => "0000000000000000",13898 => "0000000000000000",
13899 => "0000000000000000",13900 => "0000000000000000",
13901 => "0000000000000000",13902 => "0000000000000000",
13903 => "0000000000000000",13904 => "0000000000000000",
13905 => "0000000000000000",13906 => "0000000000000000",
13907 => "0000000000000000",13908 => "0000000000000000",
13909 => "0000000000000000",13910 => "0000000000000000",
13911 => "0000000000000000",13912 => "0000000000000000",
13913 => "0000000000000000",13914 => "0000000000000000",
13915 => "0000000000000000",13916 => "0000000000000000",
13917 => "0000000000000000",13918 => "0000000000000000",
13919 => "0000000000000000",13920 => "0000000000000000",
13921 => "0000000000000000",13922 => "0000000000000000",
13923 => "0000000000000000",13924 => "0000000000000000",
13925 => "0000000000000000",13926 => "0000000000000000",
13927 => "0000000000000000",13928 => "0000000000000000",
13929 => "0000000000000000",13930 => "0000000000000000",
13931 => "0000000000000000",13932 => "0000000000000000",
13933 => "0000000000000000",13934 => "0000000000000000",
13935 => "0000000000000000",13936 => "0000000000000000",
13937 => "0000000000000000",13938 => "0000000000000000",
13939 => "0000000000000000",13940 => "0000000000000000",
13941 => "0000000000000000",13942 => "0000000000000000",
13943 => "0000000000000000",13944 => "0000000000000000",
13945 => "0000000000000000",13946 => "0000000000000000",
13947 => "0000000000000000",13948 => "0000000000000000",
13949 => "0000000000000000",13950 => "0000000000000000",
13951 => "0000000000000000",13952 => "0000000000000000",
13953 => "0000000000000000",13954 => "0000000000000000",
13955 => "0000000000000000",13956 => "0000000000000000",
13957 => "0000000000000000",13958 => "0000000000000000",
13959 => "0000000000000000",13960 => "0000000000000000",
13961 => "0000000000000000",13962 => "0000000000000000",
13963 => "0000000000000000",13964 => "0000000000000000",
13965 => "0000000000000000",13966 => "0000000000000000",
13967 => "0000000000000000",13968 => "0000000000000000",
13969 => "0000000000000000",13970 => "0000000000000000",
13971 => "0000000000000000",13972 => "0000000000000000",
13973 => "0000000000000000",13974 => "0000000000000000",
13975 => "0000000000000000",13976 => "0000000000000000",
13977 => "0000000000000000",13978 => "0000000000000000",
13979 => "0000000000000000",13980 => "0000000000000000",
13981 => "0000000000000000",13982 => "0000000000000000",
13983 => "0000000000000000",13984 => "0000000000000000",
13985 => "0000000000000000",13986 => "0000000000000000",
13987 => "0000000000000000",13988 => "0000000000000000",
13989 => "0000000000000000",13990 => "0000000000000000",
13991 => "0000000000000000",13992 => "0000000000000000",
13993 => "0000000000000000",13994 => "0000000000000000",
13995 => "0000000000000000",13996 => "0000000000000000",
13997 => "0000000000000000",13998 => "0000000000000000",
13999 => "0000000000000000",14000 => "0000000000000000",
14001 => "0000000000000000",14002 => "0000000000000000",
14003 => "0000000000000000",14004 => "0000000000000000",
14005 => "0000000000000000",14006 => "0000000000000000",
14007 => "0000000000000000",14008 => "0000000000000000",
14009 => "0000000000000000",14010 => "0000000000000000",
14011 => "0000000000000000",14012 => "0000000000000000",
14013 => "0000000000000000",14014 => "0000000000000000",
14015 => "0000000000000000",14016 => "0000000000000000",
14017 => "0000000000000000",14018 => "0000000000000000",
14019 => "0000000000000000",14020 => "0000000000000000",
14021 => "0000000000000000",14022 => "0000000000000000",
14023 => "0000000000000000",14024 => "0000000000000000",
14025 => "0000000000000000",14026 => "0000000000000000",
14027 => "0000000000000000",14028 => "0000000000000000",
14029 => "0000000000000000",14030 => "0000000000000000",
14031 => "0000000000000000",14032 => "0000000000000000",
14033 => "0000000000000000",14034 => "0000000000000000",
14035 => "0000000000000000",14036 => "0000000000000000",
14037 => "0000000000000000",14038 => "0000000000000000",
14039 => "0000000000000000",14040 => "0000000000000000",
14041 => "0000000000000000",14042 => "0000000000000000",
14043 => "0000000000000000",14044 => "0000000000000000",
14045 => "0000000000000000",14046 => "0000000000000000",
14047 => "0000000000000000",14048 => "0000000000000000",
14049 => "0000000000000000",14050 => "0000000000000000",
14051 => "0000000000000000",14052 => "0000000000000000",
14053 => "0000000000000000",14054 => "0000000000000000",
14055 => "0000000000000000",14056 => "0000000000000000",
14057 => "0000000000000000",14058 => "0000000000000000",
14059 => "0000000000000000",14060 => "0000000000000000",
14061 => "0000000000000000",14062 => "0000000000000000",
14063 => "0000000000000000",14064 => "0000000000000000",
14065 => "0000000000000000",14066 => "0000000000000000",
14067 => "0000000000000000",14068 => "0000000000000000",
14069 => "0000000000000000",14070 => "0000000000000000",
14071 => "0000000000000000",14072 => "0000000000000000",
14073 => "0000000000000000",14074 => "0000000000000000",
14075 => "0000000000000000",14076 => "0000000000000000",
14077 => "0000000000000000",14078 => "0000000000000000",
14079 => "0000000000000000",14080 => "0000000000000000",
14081 => "0000000000000000",14082 => "0000000000000000",
14083 => "0000000000000000",14084 => "0000000000000000",
14085 => "0000000000000000",14086 => "0000000000000000",
14087 => "0000000000000000",14088 => "0000000000000000",
14089 => "0000000000000000",14090 => "0000000000000000",
14091 => "0000000000000000",14092 => "0000000000000000",
14093 => "0000000000000000",14094 => "0000000000000000",
14095 => "0000000000000000",14096 => "0000000000000000",
14097 => "0000000000000000",14098 => "0000000000000000",
14099 => "0000000000000000",14100 => "0000000000000000",
14101 => "0000000000000000",14102 => "0000000000000000",
14103 => "0000000000000000",14104 => "0000000000000000",
14105 => "0000000000000000",14106 => "0000000000000000",
14107 => "0000000000000000",14108 => "0000000000000000",
14109 => "0000000000000000",14110 => "0000000000000000",
14111 => "0000000000000000",14112 => "0000000000000000",
14113 => "0000000000000000",14114 => "0000000000000000",
14115 => "0000000000000000",14116 => "0000000000000000",
14117 => "0000000000000000",14118 => "0000000000000000",
14119 => "0000000000000000",14120 => "0000000000000000",
14121 => "0000000000000000",14122 => "0000000000000000",
14123 => "0000000000000000",14124 => "0000000000000000",
14125 => "0000000000000000",14126 => "0000000000000000",
14127 => "0000000000000000",14128 => "0000000000000000",
14129 => "0000000000000000",14130 => "0000000000000000",
14131 => "0000000000000000",14132 => "0000000000000000",
14133 => "0000000000000000",14134 => "0000000000000000",
14135 => "0000000000000000",14136 => "0000000000000000",
14137 => "0000000000000000",14138 => "0000000000000000",
14139 => "0000000000000000",14140 => "0000000000000000",
14141 => "0000000000000000",14142 => "0000000000000000",
14143 => "0000000000000000",14144 => "0000000000000000",
14145 => "0000000000000000",14146 => "0000000000000000",
14147 => "0000000000000000",14148 => "0000000000000000",
14149 => "0000000000000000",14150 => "0000000000000000",
14151 => "0000000000000000",14152 => "0000000000000000",
14153 => "0000000000000000",14154 => "0000000000000000",
14155 => "0000000000000000",14156 => "0000000000000000",
14157 => "0000000000000000",14158 => "0000000000000000",
14159 => "0000000000000000",14160 => "0000000000000000",
14161 => "0000000000000000",14162 => "0000000000000000",
14163 => "0000000000000000",14164 => "0000000000000000",
14165 => "0000000000000000",14166 => "0000000000000000",
14167 => "0000000000000000",14168 => "0000000000000000",
14169 => "0000000000000000",14170 => "0000000000000000",
14171 => "0000000000000000",14172 => "0000000000000000",
14173 => "0000000000000000",14174 => "0000000000000000",
14175 => "0000000000000000",14176 => "0000000000000000",
14177 => "0000000000000000",14178 => "0000000000000000",
14179 => "0000000000000000",14180 => "0000000000000000",
14181 => "0000000000000000",14182 => "0000000000000000",
14183 => "0000000000000000",14184 => "0000000000000000",
14185 => "0000000000000000",14186 => "0000000000000000",
14187 => "0000000000000000",14188 => "0000000000000000",
14189 => "0000000000000000",14190 => "0000000000000000",
14191 => "0000000000000000",14192 => "0000000000000000",
14193 => "0000000000000000",14194 => "0000000000000000",
14195 => "0000000000000000",14196 => "0000000000000000",
14197 => "0000000000000000",14198 => "0000000000000000",
14199 => "0000000000000000",14200 => "0000000000000000",
14201 => "0000000000000000",14202 => "0000000000000000",
14203 => "0000000000000000",14204 => "0000000000000000",
14205 => "0000000000000000",14206 => "0000000000000000",
14207 => "0000000000000000",14208 => "0000000000000000",
14209 => "0000000000000000",14210 => "0000000000000000",
14211 => "0000000000000000",14212 => "0000000000000000",
14213 => "0000000000000000",14214 => "0000000000000000",
14215 => "0000000000000000",14216 => "0000000000000000",
14217 => "0000000000000000",14218 => "0000000000000000",
14219 => "0000000000000000",14220 => "0000000000000000",
14221 => "0000000000000000",14222 => "0000000000000000",
14223 => "0000000000000000",14224 => "0000000000000000",
14225 => "0000000000000000",14226 => "0000000000000000",
14227 => "0000000000000000",14228 => "0000000000000000",
14229 => "0000000000000000",14230 => "0000000000000000",
14231 => "0000000000000000",14232 => "0000000000000000",
14233 => "0000000000000000",14234 => "0000000000000000",
14235 => "0000000000000000",14236 => "0000000000000000",
14237 => "0000000000000000",14238 => "0000000000000000",
14239 => "0000000000000000",14240 => "0000000000000000",
14241 => "0000000000000000",14242 => "0000000000000000",
14243 => "0000000000000000",14244 => "0000000000000000",
14245 => "0000000000000000",14246 => "0000000000000000",
14247 => "0000000000000000",14248 => "0000000000000000",
14249 => "0000000000000000",14250 => "0000000000000000",
14251 => "0000000000000000",14252 => "0000000000000000",
14253 => "0000000000000000",14254 => "0000000000000000",
14255 => "0000000000000000",14256 => "0000000000000000",
14257 => "0000000000000000",14258 => "0000000000000000",
14259 => "0000000000000000",14260 => "0000000000000000",
14261 => "0000000000000000",14262 => "0000000000000000",
14263 => "0000000000000000",14264 => "0000000000000000",
14265 => "0000000000000000",14266 => "0000000000000000",
14267 => "0000000000000000",14268 => "0000000000000000",
14269 => "0000000000000000",14270 => "0000000000000000",
14271 => "0000000000000000",14272 => "0000000000000000",
14273 => "0000000000000000",14274 => "0000000000000000",
14275 => "0000000000000000",14276 => "0000000000000000",
14277 => "0000000000000000",14278 => "0000000000000000",
14279 => "0000000000000000",14280 => "0000000000000000",
14281 => "0000000000000000",14282 => "0000000000000000",
14283 => "0000000000000000",14284 => "0000000000000000",
14285 => "0000000000000000",14286 => "0000000000000000",
14287 => "0000000000000000",14288 => "0000000000000000",
14289 => "0000000000000000",14290 => "0000000000000000",
14291 => "0000000000000000",14292 => "0000000000000000",
14293 => "0000000000000000",14294 => "0000000000000000",
14295 => "0000000000000000",14296 => "0000000000000000",
14297 => "0000000000000000",14298 => "0000000000000000",
14299 => "0000000000000000",14300 => "0000000000000000",
14301 => "0000000000000000",14302 => "0000000000000000",
14303 => "0000000000000000",14304 => "0000000000000000",
14305 => "0000000000000000",14306 => "0000000000000000",
14307 => "0000000000000000",14308 => "0000000000000000",
14309 => "0000000000000000",14310 => "0000000000000000",
14311 => "0000000000000000",14312 => "0000000000000000",
14313 => "0000000000000000",14314 => "0000000000000000",
14315 => "0000000000000000",14316 => "0000000000000000",
14317 => "0000000000000000",14318 => "0000000000000000",
14319 => "0000000000000000",14320 => "0000000000000000",
14321 => "0000000000000000",14322 => "0000000000000000",
14323 => "0000000000000000",14324 => "0000000000000000",
14325 => "0000000000000000",14326 => "0000000000000000",
14327 => "0000000000000000",14328 => "0000000000000000",
14329 => "0000000000000000",14330 => "0000000000000000",
14331 => "0000000000000000",14332 => "0000000000000000",
14333 => "0000000000000000",14334 => "0000000000000000",
14335 => "0000000000000000",14336 => "0000000000000000",
14337 => "0000000000000000",14338 => "0000000000000000",
14339 => "0000000000000000",14340 => "0000000000000000",
14341 => "0000000000000000",14342 => "0000000000000000",
14343 => "0000000000000000",14344 => "0000000000000000",
14345 => "0000000000000000",14346 => "0000000000000000",
14347 => "0000000000000000",14348 => "0000000000000000",
14349 => "0000000000000000",14350 => "0000000000000000",
14351 => "0000000000000000",14352 => "0000000000000000",
14353 => "0000000000000000",14354 => "0000000000000000",
14355 => "0000000000000000",14356 => "0000000000000000",
14357 => "0000000000000000",14358 => "0000000000000000",
14359 => "0000000000000000",14360 => "0000000000000000",
14361 => "0000000000000000",14362 => "0000000000000000",
14363 => "0000000000000000",14364 => "0000000000000000",
14365 => "0000000000000000",14366 => "0000000000000000",
14367 => "0000000000000000",14368 => "0000000000000000",
14369 => "0000000000000000",14370 => "0000000000000000",
14371 => "0000000000000000",14372 => "0000000000000000",
14373 => "0000000000000000",14374 => "0000000000000000",
14375 => "0000000000000000",14376 => "0000000000000000",
14377 => "0000000000000000",14378 => "0000000000000000",
14379 => "0000000000000000",14380 => "0000000000000000",
14381 => "0000000000000000",14382 => "0000000000000000",
14383 => "0000000000000000",14384 => "0000000000000000",
14385 => "0000000000000000",14386 => "0000000000000000",
14387 => "0000000000000000",14388 => "0000000000000000",
14389 => "0000000000000000",14390 => "0000000000000000",
14391 => "0000000000000000",14392 => "0000000000000000",
14393 => "0000000000000000",14394 => "0000000000000000",
14395 => "0000000000000000",14396 => "0000000000000000",
14397 => "0000000000000000",14398 => "0000000000000000",
14399 => "0000000000000000",14400 => "0000000000000000",
14401 => "0000000000000000",14402 => "0000000000000000",
14403 => "0000000000000000",14404 => "0000000000000000",
14405 => "0000000000000000",14406 => "0000000000000000",
14407 => "0000000000000000",14408 => "0000000000000000",
14409 => "0000000000000000",14410 => "0000000000000000",
14411 => "0000000000000000",14412 => "0000000000000000",
14413 => "0000000000000000",14414 => "0000000000000000",
14415 => "0000000000000000",14416 => "0000000000000000",
14417 => "0000000000000000",14418 => "0000000000000000",
14419 => "0000000000000000",14420 => "0000000000000000",
14421 => "0000000000000000",14422 => "0000000000000000",
14423 => "0000000000000000",14424 => "0000000000000000",
14425 => "0000000000000000",14426 => "0000000000000000",
14427 => "0000000000000000",14428 => "0000000000000000",
14429 => "0000000000000000",14430 => "0000000000000000",
14431 => "0000000000000000",14432 => "0000000000000000",
14433 => "0000000000000000",14434 => "0000000000000000",
14435 => "0000000000000000",14436 => "0000000000000000",
14437 => "0000000000000000",14438 => "0000000000000000",
14439 => "0000000000000000",14440 => "0000000000000000",
14441 => "0000000000000000",14442 => "0000000000000000",
14443 => "0000000000000000",14444 => "0000000000000000",
14445 => "0000000000000000",14446 => "0000000000000000",
14447 => "0000000000000000",14448 => "0000000000000000",
14449 => "0000000000000000",14450 => "0000000000000000",
14451 => "0000000000000000",14452 => "0000000000000000",
14453 => "0000000000000000",14454 => "0000000000000000",
14455 => "0000000000000000",14456 => "0000000000000000",
14457 => "0000000000000000",14458 => "0000000000000000",
14459 => "0000000000000000",14460 => "0000000000000000",
14461 => "0000000000000000",14462 => "0000000000000000",
14463 => "0000000000000000",14464 => "0000000000000000",
14465 => "0000000000000000",14466 => "0000000000000000",
14467 => "0000000000000000",14468 => "0000000000000000",
14469 => "0000000000000000",14470 => "0000000000000000",
14471 => "0000000000000000",14472 => "0000000000000000",
14473 => "0000000000000000",14474 => "0000000000000000",
14475 => "0000000000000000",14476 => "0000000000000000",
14477 => "0000000000000000",14478 => "0000000000000000",
14479 => "0000000000000000",14480 => "0000000000000000",
14481 => "0000000000000000",14482 => "0000000000000000",
14483 => "0000000000000000",14484 => "0000000000000000",
14485 => "0000000000000000",14486 => "0000000000000000",
14487 => "0000000000000000",14488 => "0000000000000000",
14489 => "0000000000000000",14490 => "0000000000000000",
14491 => "0000000000000000",14492 => "0000000000000000",
14493 => "0000000000000000",14494 => "0000000000000000",
14495 => "0000000000000000",14496 => "0000000000000000",
14497 => "0000000000000000",14498 => "0000000000000000",
14499 => "0000000000000000",14500 => "0000000000000000",
14501 => "0000000000000000",14502 => "0000000000000000",
14503 => "0000000000000000",14504 => "0000000000000000",
14505 => "0000000000000000",14506 => "0000000000000000",
14507 => "0000000000000000",14508 => "0000000000000000",
14509 => "0000000000000000",14510 => "0000000000000000",
14511 => "0000000000000000",14512 => "0000000000000000",
14513 => "0000000000000000",14514 => "0000000000000000",
14515 => "0000000000000000",14516 => "0000000000000000",
14517 => "0000000000000000",14518 => "0000000000000000",
14519 => "0000000000000000",14520 => "0000000000000000",
14521 => "0000000000000000",14522 => "0000000000000000",
14523 => "0000000000000000",14524 => "0000000000000000",
14525 => "0000000000000000",14526 => "0000000000000000",
14527 => "0000000000000000",14528 => "0000000000000000",
14529 => "0000000000000000",14530 => "0000000000000000",
14531 => "0000000000000000",14532 => "0000000000000000",
14533 => "0000000000000000",14534 => "0000000000000000",
14535 => "0000000000000000",14536 => "0000000000000000",
14537 => "0000000000000000",14538 => "0000000000000000",
14539 => "0000000000000000",14540 => "0000000000000000",
14541 => "0000000000000000",14542 => "0000000000000000",
14543 => "0000000000000000",14544 => "0000000000000000",
14545 => "0000000000000000",14546 => "0000000000000000",
14547 => "0000000000000000",14548 => "0000000000000000",
14549 => "0000000000000000",14550 => "0000000000000000",
14551 => "0000000000000000",14552 => "0000000000000000",
14553 => "0000000000000000",14554 => "0000000000000000",
14555 => "0000000000000000",14556 => "0000000000000000",
14557 => "0000000000000000",14558 => "0000000000000000",
14559 => "0000000000000000",14560 => "0000000000000000",
14561 => "0000000000000000",14562 => "0000000000000000",
14563 => "0000000000000000",14564 => "0000000000000000",
14565 => "0000000000000000",14566 => "0000000000000000",
14567 => "0000000000000000",14568 => "0000000000000000",
14569 => "0000000000000000",14570 => "0000000000000000",
14571 => "0000000000000000",14572 => "0000000000000000",
14573 => "0000000000000000",14574 => "0000000000000000",
14575 => "0000000000000000",14576 => "0000000000000000",
14577 => "0000000000000000",14578 => "0000000000000000",
14579 => "0000000000000000",14580 => "0000000000000000",
14581 => "0000000000000000",14582 => "0000000000000000",
14583 => "0000000000000000",14584 => "0000000000000000",
14585 => "0000000000000000",14586 => "0000000000000000",
14587 => "0000000000000000",14588 => "0000000000000000",
14589 => "0000000000000000",14590 => "0000000000000000",
14591 => "0000000000000000",14592 => "0000000000000000",
14593 => "0000000000000000",14594 => "0000000000000000",
14595 => "0000000000000000",14596 => "0000000000000000",
14597 => "0000000000000000",14598 => "0000000000000000",
14599 => "0000000000000000",14600 => "0000000000000000",
14601 => "0000000000000000",14602 => "0000000000000000",
14603 => "0000000000000000",14604 => "0000000000000000",
14605 => "0000000000000000",14606 => "0000000000000000",
14607 => "0000000000000000",14608 => "0000000000000000",
14609 => "0000000000000000",14610 => "0000000000000000",
14611 => "0000000000000000",14612 => "0000000000000000",
14613 => "0000000000000000",14614 => "0000000000000000",
14615 => "0000000000000000",14616 => "0000000000000000",
14617 => "0000000000000000",14618 => "0000000000000000",
14619 => "0000000000000000",14620 => "0000000000000000",
14621 => "0000000000000000",14622 => "0000000000000000",
14623 => "0000000000000000",14624 => "0000000000000000",
14625 => "0000000000000000",14626 => "0000000000000000",
14627 => "0000000000000000",14628 => "0000000000000000",
14629 => "0000000000000000",14630 => "0000000000000000",
14631 => "0000000000000000",14632 => "0000000000000000",
14633 => "0000000000000000",14634 => "0000000000000000",
14635 => "0000000000000000",14636 => "0000000000000000",
14637 => "0000000000000000",14638 => "0000000000000000",
14639 => "0000000000000000",14640 => "0000000000000000",
14641 => "0000000000000000",14642 => "0000000000000000",
14643 => "0000000000000000",14644 => "0000000000000000",
14645 => "0000000000000000",14646 => "0000000000000000",
14647 => "0000000000000000",14648 => "0000000000000000",
14649 => "0000000000000000",14650 => "0000000000000000",
14651 => "0000000000000000",14652 => "0000000000000000",
14653 => "0000000000000000",14654 => "0000000000000000",
14655 => "0000000000000000",14656 => "0000000000000000",
14657 => "0000000000000000",14658 => "0000000000000000",
14659 => "0000000000000000",14660 => "0000000000000000",
14661 => "0000000000000000",14662 => "0000000000000000",
14663 => "0000000000000000",14664 => "0000000000000000",
14665 => "0000000000000000",14666 => "0000000000000000",
14667 => "0000000000000000",14668 => "0000000000000000",
14669 => "0000000000000000",14670 => "0000000000000000",
14671 => "0000000000000000",14672 => "0000000000000000",
14673 => "0000000000000000",14674 => "0000000000000000",
14675 => "0000000000000000",14676 => "0000000000000000",
14677 => "0000000000000000",14678 => "0000000000000000",
14679 => "0000000000000000",14680 => "0000000000000000",
14681 => "0000000000000000",14682 => "0000000000000000",
14683 => "0000000000000000",14684 => "0000000000000000",
14685 => "0000000000000000",14686 => "0000000000000000",
14687 => "0000000000000000",14688 => "0000000000000000",
14689 => "0000000000000000",14690 => "0000000000000000",
14691 => "0000000000000000",14692 => "0000000000000000",
14693 => "0000000000000000",14694 => "0000000000000000",
14695 => "0000000000000000",14696 => "0000000000000000",
14697 => "0000000000000000",14698 => "0000000000000000",
14699 => "0000000000000000",14700 => "0000000000000000",
14701 => "0000000000000000",14702 => "0000000000000000",
14703 => "0000000000000000",14704 => "0000000000000000",
14705 => "0000000000000000",14706 => "0000000000000000",
14707 => "0000000000000000",14708 => "0000000000000000",
14709 => "0000000000000000",14710 => "0000000000000000",
14711 => "0000000000000000",14712 => "0000000000000000",
14713 => "0000000000000000",14714 => "0000000000000000",
14715 => "0000000000000000",14716 => "0000000000000000",
14717 => "0000000000000000",14718 => "0000000000000000",
14719 => "0000000000000000",14720 => "0000000000000000",
14721 => "0000000000000000",14722 => "0000000000000000",
14723 => "0000000000000000",14724 => "0000000000000000",
14725 => "0000000000000000",14726 => "0000000000000000",
14727 => "0000000000000000",14728 => "0000000000000000",
14729 => "0000000000000000",14730 => "0000000000000000",
14731 => "0000000000000000",14732 => "0000000000000000",
14733 => "0000000000000000",14734 => "0000000000000000",
14735 => "0000000000000000",14736 => "0000000000000000",
14737 => "0000000000000000",14738 => "0000000000000000",
14739 => "0000000000000000",14740 => "0000000000000000",
14741 => "0000000000000000",14742 => "0000000000000000",
14743 => "0000000000000000",14744 => "0000000000000000",
14745 => "0000000000000000",14746 => "0000000000000000",
14747 => "0000000000000000",14748 => "0000000000000000",
14749 => "0000000000000000",14750 => "0000000000000000",
14751 => "0000000000000000",14752 => "0000000000000000",
14753 => "0000000000000000",14754 => "0000000000000000",
14755 => "0000000000000000",14756 => "0000000000000000",
14757 => "0000000000000000",14758 => "0000000000000000",
14759 => "0000000000000000",14760 => "0000000000000000",
14761 => "0000000000000000",14762 => "0000000000000000",
14763 => "0000000000000000",14764 => "0000000000000000",
14765 => "0000000000000000",14766 => "0000000000000000",
14767 => "0000000000000000",14768 => "0000000000000000",
14769 => "0000000000000000",14770 => "0000000000000000",
14771 => "0000000000000000",14772 => "0000000000000000",
14773 => "0000000000000000",14774 => "0000000000000000",
14775 => "0000000000000000",14776 => "0000000000000000",
14777 => "0000000000000000",14778 => "0000000000000000",
14779 => "0000000000000000",14780 => "0000000000000000",
14781 => "0000000000000000",14782 => "0000000000000000",
14783 => "0000000000000000",14784 => "0000000000000000",
14785 => "0000000000000000",14786 => "0000000000000000",
14787 => "0000000000000000",14788 => "0000000000000000",
14789 => "0000000000000000",14790 => "0000000000000000",
14791 => "0000000000000000",14792 => "0000000000000000",
14793 => "0000000000000000",14794 => "0000000000000000",
14795 => "0000000000000000",14796 => "0000000000000000",
14797 => "0000000000000000",14798 => "0000000000000000",
14799 => "0000000000000000",14800 => "0000000000000000",
14801 => "0000000000000000",14802 => "0000000000000000",
14803 => "0000000000000000",14804 => "0000000000000000",
14805 => "0000000000000000",14806 => "0000000000000000",
14807 => "0000000000000000",14808 => "0000000000000000",
14809 => "0000000000000000",14810 => "0000000000000000",
14811 => "0000000000000000",14812 => "0000000000000000",
14813 => "0000000000000000",14814 => "0000000000000000",
14815 => "0000000000000000",14816 => "0000000000000000",
14817 => "0000000000000000",14818 => "0000000000000000",
14819 => "0000000000000000",14820 => "0000000000000000",
14821 => "0000000000000000",14822 => "0000000000000000",
14823 => "0000000000000000",14824 => "0000000000000000",
14825 => "0000000000000000",14826 => "0000000000000000",
14827 => "0000000000000000",14828 => "0000000000000000",
14829 => "0000000000000000",14830 => "0000000000000000",
14831 => "0000000000000000",14832 => "0000000000000000",
14833 => "0000000000000000",14834 => "0000000000000000",
14835 => "0000000000000000",14836 => "0000000000000000",
14837 => "0000000000000000",14838 => "0000000000000000",
14839 => "0000000000000000",14840 => "0000000000000000",
14841 => "0000000000000000",14842 => "0000000000000000",
14843 => "0000000000000000",14844 => "0000000000000000",
14845 => "0000000000000000",14846 => "0000000000000000",
14847 => "0000000000000000",14848 => "0000000000000000",
14849 => "0000000000000000",14850 => "0000000000000000",
14851 => "0000000000000000",14852 => "0000000000000000",
14853 => "0000000000000000",14854 => "0000000000000000",
14855 => "0000000000000000",14856 => "0000000000000000",
14857 => "0000000000000000",14858 => "0000000000000000",
14859 => "0000000000000000",14860 => "0000000000000000",
14861 => "0000000000000000",14862 => "0000000000000000",
14863 => "0000000000000000",14864 => "0000000000000000",
14865 => "0000000000000000",14866 => "0000000000000000",
14867 => "0000000000000000",14868 => "0000000000000000",
14869 => "0000000000000000",14870 => "0000000000000000",
14871 => "0000000000000000",14872 => "0000000000000000",
14873 => "0000000000000000",14874 => "0000000000000000",
14875 => "0000000000000000",14876 => "0000000000000000",
14877 => "0000000000000000",14878 => "0000000000000000",
14879 => "0000000000000000",14880 => "0000000000000000",
14881 => "0000000000000000",14882 => "0000000000000000",
14883 => "0000000000000000",14884 => "0000000000000000",
14885 => "0000000000000000",14886 => "0000000000000000",
14887 => "0000000000000000",14888 => "0000000000000000",
14889 => "0000000000000000",14890 => "0000000000000000",
14891 => "0000000000000000",14892 => "0000000000000000",
14893 => "0000000000000000",14894 => "0000000000000000",
14895 => "0000000000000000",14896 => "0000000000000000",
14897 => "0000000000000000",14898 => "0000000000000000",
14899 => "0000000000000000",14900 => "0000000000000000",
14901 => "0000000000000000",14902 => "0000000000000000",
14903 => "0000000000000000",14904 => "0000000000000000",
14905 => "0000000000000000",14906 => "0000000000000000",
14907 => "0000000000000000",14908 => "0000000000000000",
14909 => "0000000000000000",14910 => "0000000000000000",
14911 => "0000000000000000",14912 => "0000000000000000",
14913 => "0000000000000000",14914 => "0000000000000000",
14915 => "0000000000000000",14916 => "0000000000000000",
14917 => "0000000000000000",14918 => "0000000000000000",
14919 => "0000000000000000",14920 => "0000000000000000",
14921 => "0000000000000000",14922 => "0000000000000000",
14923 => "0000000000000000",14924 => "0000000000000000",
14925 => "0000000000000000",14926 => "0000000000000000",
14927 => "0000000000000000",14928 => "0000000000000000",
14929 => "0000000000000000",14930 => "0000000000000000",
14931 => "0000000000000000",14932 => "0000000000000000",
14933 => "0000000000000000",14934 => "0000000000000000",
14935 => "0000000000000000",14936 => "0000000000000000",
14937 => "0000000000000000",14938 => "0000000000000000",
14939 => "0000000000000000",14940 => "0000000000000000",
14941 => "0000000000000000",14942 => "0000000000000000",
14943 => "0000000000000000",14944 => "0000000000000000",
14945 => "0000000000000000",14946 => "0000000000000000",
14947 => "0000000000000000",14948 => "0000000000000000",
14949 => "0000000000000000",14950 => "0000000000000000",
14951 => "0000000000000000",14952 => "0000000000000000",
14953 => "0000000000000000",14954 => "0000000000000000",
14955 => "0000000000000000",14956 => "0000000000000000",
14957 => "0000000000000000",14958 => "0000000000000000",
14959 => "0000000000000000",14960 => "0000000000000000",
14961 => "0000000000000000",14962 => "0000000000000000",
14963 => "0000000000000000",14964 => "0000000000000000",
14965 => "0000000000000000",14966 => "0000000000000000",
14967 => "0000000000000000",14968 => "0000000000000000",
14969 => "0000000000000000",14970 => "0000000000000000",
14971 => "0000000000000000",14972 => "0000000000000000",
14973 => "0000000000000000",14974 => "0000000000000000",
14975 => "0000000000000000",14976 => "0000000000000000",
14977 => "0000000000000000",14978 => "0000000000000000",
14979 => "0000000000000000",14980 => "0000000000000000",
14981 => "0000000000000000",14982 => "0000000000000000",
14983 => "0000000000000000",14984 => "0000000000000000",
14985 => "0000000000000000",14986 => "0000000000000000",
14987 => "0000000000000000",14988 => "0000000000000000",
14989 => "0000000000000000",14990 => "0000000000000000",
14991 => "0000000000000000",14992 => "0000000000000000",
14993 => "0000000000000000",14994 => "0000000000000000",
14995 => "0000000000000000",14996 => "0000000000000000",
14997 => "0000000000000000",14998 => "0000000000000000",
14999 => "0000000000000000",15000 => "0000000000000000",
15001 => "0000000000000000",15002 => "0000000000000000",
15003 => "0000000000000000",15004 => "0000000000000000",
15005 => "0000000000000000",15006 => "0000000000000000",
15007 => "0000000000000000",15008 => "0000000000000000",
15009 => "0000000000000000",15010 => "0000000000000000",
15011 => "0000000000000000",15012 => "0000000000000000",
15013 => "0000000000000000",15014 => "0000000000000000",
15015 => "0000000000000000",15016 => "0000000000000000",
15017 => "0000000000000000",15018 => "0000000000000000",
15019 => "0000000000000000",15020 => "0000000000000000",
15021 => "0000000000000000",15022 => "0000000000000000",
15023 => "0000000000000000",15024 => "0000000000000000",
15025 => "0000000000000000",15026 => "0000000000000000",
15027 => "0000000000000000",15028 => "0000000000000000",
15029 => "0000000000000000",15030 => "0000000000000000",
15031 => "0000000000000000",15032 => "0000000000000000",
15033 => "0000000000000000",15034 => "0000000000000000",
15035 => "0000000000000000",15036 => "0000000000000000",
15037 => "0000000000000000",15038 => "0000000000000000",
15039 => "0000000000000000",15040 => "0000000000000000",
15041 => "0000000000000000",15042 => "0000000000000000",
15043 => "0000000000000000",15044 => "0000000000000000",
15045 => "0000000000000000",15046 => "0000000000000000",
15047 => "0000000000000000",15048 => "0000000000000000",
15049 => "0000000000000000",15050 => "0000000000000000",
15051 => "0000000000000000",15052 => "0000000000000000",
15053 => "0000000000000000",15054 => "0000000000000000",
15055 => "0000000000000000",15056 => "0000000000000000",
15057 => "0000000000000000",15058 => "0000000000000000",
15059 => "0000000000000000",15060 => "0000000000000000",
15061 => "0000000000000000",15062 => "0000000000000000",
15063 => "0000000000000000",15064 => "0000000000000000",
15065 => "0000000000000000",15066 => "0000000000000000",
15067 => "0000000000000000",15068 => "0000000000000000",
15069 => "0000000000000000",15070 => "0000000000000000",
15071 => "0000000000000000",15072 => "0000000000000000",
15073 => "0000000000000000",15074 => "0000000000000000",
15075 => "0000000000000000",15076 => "0000000000000000",
15077 => "0000000000000000",15078 => "0000000000000000",
15079 => "0000000000000000",15080 => "0000000000000000",
15081 => "0000000000000000",15082 => "0000000000000000",
15083 => "0000000000000000",15084 => "0000000000000000",
15085 => "0000000000000000",15086 => "0000000000000000",
15087 => "0000000000000000",15088 => "0000000000000000",
15089 => "0000000000000000",15090 => "0000000000000000",
15091 => "0000000000000000",15092 => "0000000000000000",
15093 => "0000000000000000",15094 => "0000000000000000",
15095 => "0000000000000000",15096 => "0000000000000000",
15097 => "0000000000000000",15098 => "0000000000000000",
15099 => "0000000000000000",15100 => "0000000000000000",
15101 => "0000000000000000",15102 => "0000000000000000",
15103 => "0000000000000000",15104 => "0000000000000000",
15105 => "0000000000000000",15106 => "0000000000000000",
15107 => "0000000000000000",15108 => "0000000000000000",
15109 => "0000000000000000",15110 => "0000000000000000",
15111 => "0000000000000000",15112 => "0000000000000000",
15113 => "0000000000000000",15114 => "0000000000000000",
15115 => "0000000000000000",15116 => "0000000000000000",
15117 => "0000000000000000",15118 => "0000000000000000",
15119 => "0000000000000000",15120 => "0000000000000000",
15121 => "0000000000000000",15122 => "0000000000000000",
15123 => "0000000000000000",15124 => "0000000000000000",
15125 => "0000000000000000",15126 => "0000000000000000",
15127 => "0000000000000000",15128 => "0000000000000000",
15129 => "0000000000000000",15130 => "0000000000000000",
15131 => "0000000000000000",15132 => "0000000000000000",
15133 => "0000000000000000",15134 => "0000000000000000",
15135 => "0000000000000000",15136 => "0000000000000000",
15137 => "0000000000000000",15138 => "0000000000000000",
15139 => "0000000000000000",15140 => "0000000000000000",
15141 => "0000000000000000",15142 => "0000000000000000",
15143 => "0000000000000000",15144 => "0000000000000000",
15145 => "0000000000000000",15146 => "0000000000000000",
15147 => "0000000000000000",15148 => "0000000000000000",
15149 => "0000000000000000",15150 => "0000000000000000",
15151 => "0000000000000000",15152 => "0000000000000000",
15153 => "0000000000000000",15154 => "0000000000000000",
15155 => "0000000000000000",15156 => "0000000000000000",
15157 => "0000000000000000",15158 => "0000000000000000",
15159 => "0000000000000000",15160 => "0000000000000000",
15161 => "0000000000000000",15162 => "0000000000000000",
15163 => "0000000000000000",15164 => "0000000000000000",
15165 => "0000000000000000",15166 => "0000000000000000",
15167 => "0000000000000000",15168 => "0000000000000000",
15169 => "0000000000000000",15170 => "0000000000000000",
15171 => "0000000000000000",15172 => "0000000000000000",
15173 => "0000000000000000",15174 => "0000000000000000",
15175 => "0000000000000000",15176 => "0000000000000000",
15177 => "0000000000000000",15178 => "0000000000000000",
15179 => "0000000000000000",15180 => "0000000000000000",
15181 => "0000000000000000",15182 => "0000000000000000",
15183 => "0000000000000000",15184 => "0000000000000000",
15185 => "0000000000000000",15186 => "0000000000000000",
15187 => "0000000000000000",15188 => "0000000000000000",
15189 => "0000000000000000",15190 => "0000000000000000",
15191 => "0000000000000000",15192 => "0000000000000000",
15193 => "0000000000000000",15194 => "0000000000000000",
15195 => "0000000000000000",15196 => "0000000000000000",
15197 => "0000000000000000",15198 => "0000000000000000",
15199 => "0000000000000000",15200 => "0000000000000000",
15201 => "0000000000000000",15202 => "0000000000000000",
15203 => "0000000000000000",15204 => "0000000000000000",
15205 => "0000000000000000",15206 => "0000000000000000",
15207 => "0000000000000000",15208 => "0000000000000000",
15209 => "0000000000000000",15210 => "0000000000000000",
15211 => "0000000000000000",15212 => "0000000000000000",
15213 => "0000000000000000",15214 => "0000000000000000",
15215 => "0000000000000000",15216 => "0000000000000000",
15217 => "0000000000000000",15218 => "0000000000000000",
15219 => "0000000000000000",15220 => "0000000000000000",
15221 => "0000000000000000",15222 => "0000000000000000",
15223 => "0000000000000000",15224 => "0000000000000000",
15225 => "0000000000000000",15226 => "0000000000000000",
15227 => "0000000000000000",15228 => "0000000000000000",
15229 => "0000000000000000",15230 => "0000000000000000",
15231 => "0000000000000000",15232 => "0000000000000000",
15233 => "0000000000000000",15234 => "0000000000000000",
15235 => "0000000000000000",15236 => "0000000000000000",
15237 => "0000000000000000",15238 => "0000000000000000",
15239 => "0000000000000000",15240 => "0000000000000000",
15241 => "0000000000000000",15242 => "0000000000000000",
15243 => "0000000000000000",15244 => "0000000000000000",
15245 => "0000000000000000",15246 => "0000000000000000",
15247 => "0000000000000000",15248 => "0000000000000000",
15249 => "0000000000000000",15250 => "0000000000000000",
15251 => "0000000000000000",15252 => "0000000000000000",
15253 => "0000000000000000",15254 => "0000000000000000",
15255 => "0000000000000000",15256 => "0000000000000000",
15257 => "0000000000000000",15258 => "0000000000000000",
15259 => "0000000000000000",15260 => "0000000000000000",
15261 => "0000000000000000",15262 => "0000000000000000",
15263 => "0000000000000000",15264 => "0000000000000000",
15265 => "0000000000000000",15266 => "0000000000000000",
15267 => "0000000000000000",15268 => "0000000000000000",
15269 => "0000000000000000",15270 => "0000000000000000",
15271 => "0000000000000000",15272 => "0000000000000000",
15273 => "0000000000000000",15274 => "0000000000000000",
15275 => "0000000000000000",15276 => "0000000000000000",
15277 => "0000000000000000",15278 => "0000000000000000",
15279 => "0000000000000000",15280 => "0000000000000000",
15281 => "0000000000000000",15282 => "0000000000000000",
15283 => "0000000000000000",15284 => "0000000000000000",
15285 => "0000000000000000",15286 => "0000000000000000",
15287 => "0000000000000000",15288 => "0000000000000000",
15289 => "0000000000000000",15290 => "0000000000000000",
15291 => "0000000000000000",15292 => "0000000000000000",
15293 => "0000000000000000",15294 => "0000000000000000",
15295 => "0000000000000000",15296 => "0000000000000000",
15297 => "0000000000000000",15298 => "0000000000000000",
15299 => "0000000000000000",15300 => "0000000000000000",
15301 => "0000000000000000",15302 => "0000000000000000",
15303 => "0000000000000000",15304 => "0000000000000000",
15305 => "0000000000000000",15306 => "0000000000000000",
15307 => "0000000000000000",15308 => "0000000000000000",
15309 => "0000000000000000",15310 => "0000000000000000",
15311 => "0000000000000000",15312 => "0000000000000000",
15313 => "0000000000000000",15314 => "0000000000000000",
15315 => "0000000000000000",15316 => "0000000000000000",
15317 => "0000000000000000",15318 => "0000000000000000",
15319 => "0000000000000000",15320 => "0000000000000000",
15321 => "0000000000000000",15322 => "0000000000000000",
15323 => "0000000000000000",15324 => "0000000000000000",
15325 => "0000000000000000",15326 => "0000000000000000",
15327 => "0000000000000000",15328 => "0000000000000000",
15329 => "0000000000000000",15330 => "0000000000000000",
15331 => "0000000000000000",15332 => "0000000000000000",
15333 => "0000000000000000",15334 => "0000000000000000",
15335 => "0000000000000000",15336 => "0000000000000000",
15337 => "0000000000000000",15338 => "0000000000000000",
15339 => "0000000000000000",15340 => "0000000000000000",
15341 => "0000000000000000",15342 => "0000000000000000",
15343 => "0000000000000000",15344 => "0000000000000000",
15345 => "0000000000000000",15346 => "0000000000000000",
15347 => "0000000000000000",15348 => "0000000000000000",
15349 => "0000000000000000",15350 => "0000000000000000",
15351 => "0000000000000000",15352 => "0000000000000000",
15353 => "0000000000000000",15354 => "0000000000000000",
15355 => "0000000000000000",15356 => "0000000000000000",
15357 => "0000000000000000",15358 => "0000000000000000",
15359 => "0000000000000000",15360 => "0000000000000000",
15361 => "0000000000000000",15362 => "0000000000000000",
15363 => "0000000000000000",15364 => "0000000000000000",
15365 => "0000000000000000",15366 => "0000000000000000",
15367 => "0000000000000000",15368 => "0000000000000000",
15369 => "0000000000000000",15370 => "0000000000000000",
15371 => "0000000000000000",15372 => "0000000000000000",
15373 => "0000000000000000",15374 => "0000000000000000",
15375 => "0000000000000000",15376 => "0000000000000000",
15377 => "0000000000000000",15378 => "0000000000000000",
15379 => "0000000000000000",15380 => "0000000000000000",
15381 => "0000000000000000",15382 => "0000000000000000",
15383 => "0000000000000000",15384 => "0000000000000000",
15385 => "0000000000000000",15386 => "0000000000000000",
15387 => "0000000000000000",15388 => "0000000000000000",
15389 => "0000000000000000",15390 => "0000000000000000",
15391 => "0000000000000000",15392 => "0000000000000000",
15393 => "0000000000000000",15394 => "0000000000000000",
15395 => "0000000000000000",15396 => "0000000000000000",
15397 => "0000000000000000",15398 => "0000000000000000",
15399 => "0000000000000000",15400 => "0000000000000000",
15401 => "0000000000000000",15402 => "0000000000000000",
15403 => "0000000000000000",15404 => "0000000000000000",
15405 => "0000000000000000",15406 => "0000000000000000",
15407 => "0000000000000000",15408 => "0000000000000000",
15409 => "0000000000000000",15410 => "0000000000000000",
15411 => "0000000000000000",15412 => "0000000000000000",
15413 => "0000000000000000",15414 => "0000000000000000",
15415 => "0000000000000000",15416 => "0000000000000000",
15417 => "0000000000000000",15418 => "0000000000000000",
15419 => "0000000000000000",15420 => "0000000000000000",
15421 => "0000000000000000",15422 => "0000000000000000",
15423 => "0000000000000000",15424 => "0000000000000000",
15425 => "0000000000000000",15426 => "0000000000000000",
15427 => "0000000000000000",15428 => "0000000000000000",
15429 => "0000000000000000",15430 => "0000000000000000",
15431 => "0000000000000000",15432 => "0000000000000000",
15433 => "0000000000000000",15434 => "0000000000000000",
15435 => "0000000000000000",15436 => "0000000000000000",
15437 => "0000000000000000",15438 => "0000000000000000",
15439 => "0000000000000000",15440 => "0000000000000000",
15441 => "0000000000000000",15442 => "0000000000000000",
15443 => "0000000000000000",15444 => "0000000000000000",
15445 => "0000000000000000",15446 => "0000000000000000",
15447 => "0000000000000000",15448 => "0000000000000000",
15449 => "0000000000000000",15450 => "0000000000000000",
15451 => "0000000000000000",15452 => "0000000000000000",
15453 => "0000000000000000",15454 => "0000000000000000",
15455 => "0000000000000000",15456 => "0000000000000000",
15457 => "0000000000000000",15458 => "0000000000000000",
15459 => "0000000000000000",15460 => "0000000000000000",
15461 => "0000000000000000",15462 => "0000000000000000",
15463 => "0000000000000000",15464 => "0000000000000000",
15465 => "0000000000000000",15466 => "0000000000000000",
15467 => "0000000000000000",15468 => "0000000000000000",
15469 => "0000000000000000",15470 => "0000000000000000",
15471 => "0000000000000000",15472 => "0000000000000000",
15473 => "0000000000000000",15474 => "0000000000000000",
15475 => "0000000000000000",15476 => "0000000000000000",
15477 => "0000000000000000",15478 => "0000000000000000",
15479 => "0000000000000000",15480 => "0000000000000000",
15481 => "0000000000000000",15482 => "0000000000000000",
15483 => "0000000000000000",15484 => "0000000000000000",
15485 => "0000000000000000",15486 => "0000000000000000",
15487 => "0000000000000000",15488 => "0000000000000000",
15489 => "0000000000000000",15490 => "0000000000000000",
15491 => "0000000000000000",15492 => "0000000000000000",
15493 => "0000000000000000",15494 => "0000000000000000",
15495 => "0000000000000000",15496 => "0000000000000000",
15497 => "0000000000000000",15498 => "0000000000000000",
15499 => "0000000000000000",15500 => "0000000000000000",
15501 => "0000000000000000",15502 => "0000000000000000",
15503 => "0000000000000000",15504 => "0000000000000000",
15505 => "0000000000000000",15506 => "0000000000000000",
15507 => "0000000000000000",15508 => "0000000000000000",
15509 => "0000000000000000",15510 => "0000000000000000",
15511 => "0000000000000000",15512 => "0000000000000000",
15513 => "0000000000000000",15514 => "0000000000000000",
15515 => "0000000000000000",15516 => "0000000000000000",
15517 => "0000000000000000",15518 => "0000000000000000",
15519 => "0000000000000000",15520 => "0000000000000000",
15521 => "0000000000000000",15522 => "0000000000000000",
15523 => "0000000000000000",15524 => "0000000000000000",
15525 => "0000000000000000",15526 => "0000000000000000",
15527 => "0000000000000000",15528 => "0000000000000000",
15529 => "0000000000000000",15530 => "0000000000000000",
15531 => "0000000000000000",15532 => "0000000000000000",
15533 => "0000000000000000",15534 => "0000000000000000",
15535 => "0000000000000000",15536 => "0000000000000000",
15537 => "0000000000000000",15538 => "0000000000000000",
15539 => "0000000000000000",15540 => "0000000000000000",
15541 => "0000000000000000",15542 => "0000000000000000",
15543 => "0000000000000000",15544 => "0000000000000000",
15545 => "0000000000000000",15546 => "0000000000000000",
15547 => "0000000000000000",15548 => "0000000000000000",
15549 => "0000000000000000",15550 => "0000000000000000",
15551 => "0000000000000000",15552 => "0000000000000000",
15553 => "0000000000000000",15554 => "0000000000000000",
15555 => "0000000000000000",15556 => "0000000000000000",
15557 => "0000000000000000",15558 => "0000000000000000",
15559 => "0000000000000000",15560 => "0000000000000000",
15561 => "0000000000000000",15562 => "0000000000000000",
15563 => "0000000000000000",15564 => "0000000000000000",
15565 => "0000000000000000",15566 => "0000000000000000",
15567 => "0000000000000000",15568 => "0000000000000000",
15569 => "0000000000000000",15570 => "0000000000000000",
15571 => "0000000000000000",15572 => "0000000000000000",
15573 => "0000000000000000",15574 => "0000000000000000",
15575 => "0000000000000000",15576 => "0000000000000000",
15577 => "0000000000000000",15578 => "0000000000000000",
15579 => "0000000000000000",15580 => "0000000000000000",
15581 => "0000000000000000",15582 => "0000000000000000",
15583 => "0000000000000000",15584 => "0000000000000000",
15585 => "0000000000000000",15586 => "0000000000000000",
15587 => "0000000000000000",15588 => "0000000000000000",
15589 => "0000000000000000",15590 => "0000000000000000",
15591 => "0000000000000000",15592 => "0000000000000000",
15593 => "0000000000000000",15594 => "0000000000000000",
15595 => "0000000000000000",15596 => "0000000000000000",
15597 => "0000000000000000",15598 => "0000000000000000",
15599 => "0000000000000000",15600 => "0000000000000000",
15601 => "0000000000000000",15602 => "0000000000000000",
15603 => "0000000000000000",15604 => "0000000000000000",
15605 => "0000000000000000",15606 => "0000000000000000",
15607 => "0000000000000000",15608 => "0000000000000000",
15609 => "0000000000000000",15610 => "0000000000000000",
15611 => "0000000000000000",15612 => "0000000000000000",
15613 => "0000000000000000",15614 => "0000000000000000",
15615 => "0000000000000000",15616 => "0000000000000000",
15617 => "0000000000000000",15618 => "0000000000000000",
15619 => "0000000000000000",15620 => "0000000000000000",
15621 => "0000000000000000",15622 => "0000000000000000",
15623 => "0000000000000000",15624 => "0000000000000000",
15625 => "0000000000000000",15626 => "0000000000000000",
15627 => "0000000000000000",15628 => "0000000000000000",
15629 => "0000000000000000",15630 => "0000000000000000",
15631 => "0000000000000000",15632 => "0000000000000000",
15633 => "0000000000000000",15634 => "0000000000000000",
15635 => "0000000000000000",15636 => "0000000000000000",
15637 => "0000000000000000",15638 => "0000000000000000",
15639 => "0000000000000000",15640 => "0000000000000000",
15641 => "0000000000000000",15642 => "0000000000000000",
15643 => "0000000000000000",15644 => "0000000000000000",
15645 => "0000000000000000",15646 => "0000000000000000",
15647 => "0000000000000000",15648 => "0000000000000000",
15649 => "0000000000000000",15650 => "0000000000000000",
15651 => "0000000000000000",15652 => "0000000000000000",
15653 => "0000000000000000",15654 => "0000000000000000",
15655 => "0000000000000000",15656 => "0000000000000000",
15657 => "0000000000000000",15658 => "0000000000000000",
15659 => "0000000000000000",15660 => "0000000000000000",
15661 => "0000000000000000",15662 => "0000000000000000",
15663 => "0000000000000000",15664 => "0000000000000000",
15665 => "0000000000000000",15666 => "0000000000000000",
15667 => "0000000000000000",15668 => "0000000000000000",
15669 => "0000000000000000",15670 => "0000000000000000",
15671 => "0000000000000000",15672 => "0000000000000000",
15673 => "0000000000000000",15674 => "0000000000000000",
15675 => "0000000000000000",15676 => "0000000000000000",
15677 => "0000000000000000",15678 => "0000000000000000",
15679 => "0000000000000000",15680 => "0000000000000000",
15681 => "0000000000000000",15682 => "0000000000000000",
15683 => "0000000000000000",15684 => "0000000000000000",
15685 => "0000000000000000",15686 => "0000000000000000",
15687 => "0000000000000000",15688 => "0000000000000000",
15689 => "0000000000000000",15690 => "0000000000000000",
15691 => "0000000000000000",15692 => "0000000000000000",
15693 => "0000000000000000",15694 => "0000000000000000",
15695 => "0000000000000000",15696 => "0000000000000000",
15697 => "0000000000000000",15698 => "0000000000000000",
15699 => "0000000000000000",15700 => "0000000000000000",
15701 => "0000000000000000",15702 => "0000000000000000",
15703 => "0000000000000000",15704 => "0000000000000000",
15705 => "0000000000000000",15706 => "0000000000000000",
15707 => "0000000000000000",15708 => "0000000000000000",
15709 => "0000000000000000",15710 => "0000000000000000",
15711 => "0000000000000000",15712 => "0000000000000000",
15713 => "0000000000000000",15714 => "0000000000000000",
15715 => "0000000000000000",15716 => "0000000000000000",
15717 => "0000000000000000",15718 => "0000000000000000",
15719 => "0000000000000000",15720 => "0000000000000000",
15721 => "0000000000000000",15722 => "0000000000000000",
15723 => "0000000000000000",15724 => "0000000000000000",
15725 => "0000000000000000",15726 => "0000000000000000",
15727 => "0000000000000000",15728 => "0000000000000000",
15729 => "0000000000000000",15730 => "0000000000000000",
15731 => "0000000000000000",15732 => "0000000000000000",
15733 => "0000000000000000",15734 => "0000000000000000",
15735 => "0000000000000000",15736 => "0000000000000000",
15737 => "0000000000000000",15738 => "0000000000000000",
15739 => "0000000000000000",15740 => "0000000000000000",
15741 => "0000000000000000",15742 => "0000000000000000",
15743 => "0000000000000000",15744 => "0000000000000000",
15745 => "0000000000000000",15746 => "0000000000000000",
15747 => "0000000000000000",15748 => "0000000000000000",
15749 => "0000000000000000",15750 => "0000000000000000",
15751 => "0000000000000000",15752 => "0000000000000000",
15753 => "0000000000000000",15754 => "0000000000000000",
15755 => "0000000000000000",15756 => "0000000000000000",
15757 => "0000000000000000",15758 => "0000000000000000",
15759 => "0000000000000000",15760 => "0000000000000000",
15761 => "0000000000000000",15762 => "0000000000000000",
15763 => "0000000000000000",15764 => "0000000000000000",
15765 => "0000000000000000",15766 => "0000000000000000",
15767 => "0000000000000000",15768 => "0000000000000000",
15769 => "0000000000000000",15770 => "0000000000000000",
15771 => "0000000000000000",15772 => "0000000000000000",
15773 => "0000000000000000",15774 => "0000000000000000",
15775 => "0000000000000000",15776 => "0000000000000000",
15777 => "0000000000000000",15778 => "0000000000000000",
15779 => "0000000000000000",15780 => "0000000000000000",
15781 => "0000000000000000",15782 => "0000000000000000",
15783 => "0000000000000000",15784 => "0000000000000000",
15785 => "0000000000000000",15786 => "0000000000000000",
15787 => "0000000000000000",15788 => "0000000000000000",
15789 => "0000000000000000",15790 => "0000000000000000",
15791 => "0000000000000000",15792 => "0000000000000000",
15793 => "0000000000000000",15794 => "0000000000000000",
15795 => "0000000000000000",15796 => "0000000000000000",
15797 => "0000000000000000",15798 => "0000000000000000",
15799 => "0000000000000000",15800 => "0000000000000000",
15801 => "0000000000000000",15802 => "0000000000000000",
15803 => "0000000000000000",15804 => "0000000000000000",
15805 => "0000000000000000",15806 => "0000000000000000",
15807 => "0000000000000000",15808 => "0000000000000000",
15809 => "0000000000000000",15810 => "0000000000000000",
15811 => "0000000000000000",15812 => "0000000000000000",
15813 => "0000000000000000",15814 => "0000000000000000",
15815 => "0000000000000000",15816 => "0000000000000000",
15817 => "0000000000000000",15818 => "0000000000000000",
15819 => "0000000000000000",15820 => "0000000000000000",
15821 => "0000000000000000",15822 => "0000000000000000",
15823 => "0000000000000000",15824 => "0000000000000000",
15825 => "0000000000000000",15826 => "0000000000000000",
15827 => "0000000000000000",15828 => "0000000000000000",
15829 => "0000000000000000",15830 => "0000000000000000",
15831 => "0000000000000000",15832 => "0000000000000000",
15833 => "0000000000000000",15834 => "0000000000000000",
15835 => "0000000000000000",15836 => "0000000000000000",
15837 => "0000000000000000",15838 => "0000000000000000",
15839 => "0000000000000000",15840 => "0000000000000000",
15841 => "0000000000000000",15842 => "0000000000000000",
15843 => "0000000000000000",15844 => "0000000000000000",
15845 => "0000000000000000",15846 => "0000000000000000",
15847 => "0000000000000000",15848 => "0000000000000000",
15849 => "0000000000000000",15850 => "0000000000000000",
15851 => "0000000000000000",15852 => "0000000000000000",
15853 => "0000000000000000",15854 => "0000000000000000",
15855 => "0000000000000000",15856 => "0000000000000000",
15857 => "0000000000000000",15858 => "0000000000000000",
15859 => "0000000000000000",15860 => "0000000000000000",
15861 => "0000000000000000",15862 => "0000000000000000",
15863 => "0000000000000000",15864 => "0000000000000000",
15865 => "0000000000000000",15866 => "0000000000000000",
15867 => "0000000000000000",15868 => "0000000000000000",
15869 => "0000000000000000",15870 => "0000000000000000",
15871 => "0000000000000000",15872 => "0000000000000000",
15873 => "0000000000000000",15874 => "0000000000000000",
15875 => "0000000000000000",15876 => "0000000000000000",
15877 => "0000000000000000",15878 => "0000000000000000",
15879 => "0000000000000000",15880 => "0000000000000000",
15881 => "0000000000000000",15882 => "0000000000000000",
15883 => "0000000000000000",15884 => "0000000000000000",
15885 => "0000000000000000",15886 => "0000000000000000",
15887 => "0000000000000000",15888 => "0000000000000000",
15889 => "0000000000000000",15890 => "0000000000000000",
15891 => "0000000000000000",15892 => "0000000000000000",
15893 => "0000000000000000",15894 => "0000000000000000",
15895 => "0000000000000000",15896 => "0000000000000000",
15897 => "0000000000000000",15898 => "0000000000000000",
15899 => "0000000000000000",15900 => "0000000000000000",
15901 => "0000000000000000",15902 => "0000000000000000",
15903 => "0000000000000000",15904 => "0000000000000000",
15905 => "0000000000000000",15906 => "0000000000000000",
15907 => "0000000000000000",15908 => "0000000000000000",
15909 => "0000000000000000",15910 => "0000000000000000",
15911 => "0000000000000000",15912 => "0000000000000000",
15913 => "0000000000000000",15914 => "0000000000000000",
15915 => "0000000000000000",15916 => "0000000000000000",
15917 => "0000000000000000",15918 => "0000000000000000",
15919 => "0000000000000000",15920 => "0000000000000000",
15921 => "0000000000000000",15922 => "0000000000000000",
15923 => "0000000000000000",15924 => "0000000000000000",
15925 => "0000000000000000",15926 => "0000000000000000",
15927 => "0000000000000000",15928 => "0000000000000000",
15929 => "0000000000000000",15930 => "0000000000000000",
15931 => "0000000000000000",15932 => "0000000000000000",
15933 => "0000000000000000",15934 => "0000000000000000",
15935 => "0000000000000000",15936 => "0000000000000000",
15937 => "0000000000000000",15938 => "0000000000000000",
15939 => "0000000000000000",15940 => "0000000000000000",
15941 => "0000000000000000",15942 => "0000000000000000",
15943 => "0000000000000000",15944 => "0000000000000000",
15945 => "0000000000000000",15946 => "0000000000000000",
15947 => "0000000000000000",15948 => "0000000000000000",
15949 => "0000000000000000",15950 => "0000000000000000",
15951 => "0000000000000000",15952 => "0000000000000000",
15953 => "0000000000000000",15954 => "0000000000000000",
15955 => "0000000000000000",15956 => "0000000000000000",
15957 => "0000000000000000",15958 => "0000000000000000",
15959 => "0000000000000000",15960 => "0000000000000000",
15961 => "0000000000000000",15962 => "0000000000000000",
15963 => "0000000000000000",15964 => "0000000000000000",
15965 => "0000000000000000",15966 => "0000000000000000",
15967 => "0000000000000000",15968 => "0000000000000000",
15969 => "0000000000000000",15970 => "0000000000000000",
15971 => "0000000000000000",15972 => "0000000000000000",
15973 => "0000000000000000",15974 => "0000000000000000",
15975 => "0000000000000000",15976 => "0000000000000000",
15977 => "0000000000000000",15978 => "0000000000000000",
15979 => "0000000000000000",15980 => "0000000000000000",
15981 => "0000000000000000",15982 => "0000000000000000",
15983 => "0000000000000000",15984 => "0000000000000000",
15985 => "0000000000000000",15986 => "0000000000000000",
15987 => "0000000000000000",15988 => "0000000000000000",
15989 => "0000000000000000",15990 => "0000000000000000",
15991 => "0000000000000000",15992 => "0000000000000000",
15993 => "0000000000000000",15994 => "0000000000000000",
15995 => "0000000000000000",15996 => "0000000000000000",
15997 => "0000000000000000",15998 => "0000000000000000",
15999 => "0000000000000000",16000 => "0000000000000000",
16001 => "0000000000000000",16002 => "0000000000000000",
16003 => "0000000000000000",16004 => "0000000000000000",
16005 => "0000000000000000",16006 => "0000000000000000",
16007 => "0000000000000000",16008 => "0000000000000000",
16009 => "0000000000000000",16010 => "0000000000000000",
16011 => "0000000000000000",16012 => "0000000000000000",
16013 => "0000000000000000",16014 => "0000000000000000",
16015 => "0000000000000000",16016 => "0000000000000000",
16017 => "0000000000000000",16018 => "0000000000000000",
16019 => "0000000000000000",16020 => "0000000000000000",
16021 => "0000000000000000",16022 => "0000000000000000",
16023 => "0000000000000000",16024 => "0000000000000000",
16025 => "0000000000000000",16026 => "0000000000000000",
16027 => "0000000000000000",16028 => "0000000000000000",
16029 => "0000000000000000",16030 => "0000000000000000",
16031 => "0000000000000000",16032 => "0000000000000000",
16033 => "0000000000000000",16034 => "0000000000000000",
16035 => "0000000000000000",16036 => "0000000000000000",
16037 => "0000000000000000",16038 => "0000000000000000",
16039 => "0000000000000000",16040 => "0000000000000000",
16041 => "0000000000000000",16042 => "0000000000000000",
16043 => "0000000000000000",16044 => "0000000000000000",
16045 => "0000000000000000",16046 => "0000000000000000",
16047 => "0000000000000000",16048 => "0000000000000000",
16049 => "0000000000000000",16050 => "0000000000000000",
16051 => "0000000000000000",16052 => "0000000000000000",
16053 => "0000000000000000",16054 => "0000000000000000",
16055 => "0000000000000000",16056 => "0000000000000000",
16057 => "0000000000000000",16058 => "0000000000000000",
16059 => "0000000000000000",16060 => "0000000000000000",
16061 => "0000000000000000",16062 => "0000000000000000",
16063 => "0000000000000000",16064 => "0000000000000000",
16065 => "0000000000000000",16066 => "0000000000000000",
16067 => "0000000000000000",16068 => "0000000000000000",
16069 => "0000000000000000",16070 => "0000000000000000",
16071 => "0000000000000000",16072 => "0000000000000000",
16073 => "0000000000000000",16074 => "0000000000000000",
16075 => "0000000000000000",16076 => "0000000000000000",
16077 => "0000000000000000",16078 => "0000000000000000",
16079 => "0000000000000000",16080 => "0000000000000000",
16081 => "0000000000000000",16082 => "0000000000000000",
16083 => "0000000000000000",16084 => "0000000000000000",
16085 => "0000000000000000",16086 => "0000000000000000",
16087 => "0000000000000000",16088 => "0000000000000000",
16089 => "0000000000000000",16090 => "0000000000000000",
16091 => "0000000000000000",16092 => "0000000000000000",
16093 => "0000000000000000",16094 => "0000000000000000",
16095 => "0000000000000000",16096 => "0000000000000000",
16097 => "0000000000000000",16098 => "0000000000000000",
16099 => "0000000000000000",16100 => "0000000000000000",
16101 => "0000000000000000",16102 => "0000000000000000",
16103 => "0000000000000000",16104 => "0000000000000000",
16105 => "0000000000000000",16106 => "0000000000000000",
16107 => "0000000000000000",16108 => "0000000000000000",
16109 => "0000000000000000",16110 => "0000000000000000",
16111 => "0000000000000000",16112 => "0000000000000000",
16113 => "0000000000000000",16114 => "0000000000000000",
16115 => "0000000000000000",16116 => "0000000000000000",
16117 => "0000000000000000",16118 => "0000000000000000",
16119 => "0000000000000000",16120 => "0000000000000000",
16121 => "0000000000000000",16122 => "0000000000000000",
16123 => "0000000000000000",16124 => "0000000000000000",
16125 => "0000000000000000",16126 => "0000000000000000",
16127 => "0000000000000000",16128 => "0000000000000000",
16129 => "0000000000000000",16130 => "0000000000000000",
16131 => "0000000000000000",16132 => "0000000000000000",
16133 => "0000000000000000",16134 => "0000000000000000",
16135 => "0000000000000000",16136 => "0000000000000000",
16137 => "0000000000000000",16138 => "0000000000000000",
16139 => "0000000000000000",16140 => "0000000000000000",
16141 => "0000000000000000",16142 => "0000000000000000",
16143 => "0000000000000000",16144 => "0000000000000000",
16145 => "0000000000000000",16146 => "0000000000000000",
16147 => "0000000000000000",16148 => "0000000000000000",
16149 => "0000000000000000",16150 => "0000000000000000",
16151 => "0000000000000000",16152 => "0000000000000000",
16153 => "0000000000000000",16154 => "0000000000000000",
16155 => "0000000000000000",16156 => "0000000000000000",
16157 => "0000000000000000",16158 => "0000000000000000",
16159 => "0000000000000000",16160 => "0000000000000000",
16161 => "0000000000000000",16162 => "0000000000000000",
16163 => "0000000000000000",16164 => "0000000000000000",
16165 => "0000000000000000",16166 => "0000000000000000",
16167 => "0000000000000000",16168 => "0000000000000000",
16169 => "0000000000000000",16170 => "0000000000000000",
16171 => "0000000000000000",16172 => "0000000000000000",
16173 => "0000000000000000",16174 => "0000000000000000",
16175 => "0000000000000000",16176 => "0000000000000000",
16177 => "0000000000000000",16178 => "0000000000000000",
16179 => "0000000000000000",16180 => "0000000000000000",
16181 => "0000000000000000",16182 => "0000000000000000",
16183 => "0000000000000000",16184 => "0000000000000000",
16185 => "0000000000000000",16186 => "0000000000000000",
16187 => "0000000000000000",16188 => "0000000000000000",
16189 => "0000000000000000",16190 => "0000000000000000",
16191 => "0000000000000000",16192 => "0000000000000000",
16193 => "0000000000000000",16194 => "0000000000000000",
16195 => "0000000000000000",16196 => "0000000000000000",
16197 => "0000000000000000",16198 => "0000000000000000",
16199 => "0000000000000000",16200 => "0000000000000000",
16201 => "0000000000000000",16202 => "0000000000000000",
16203 => "0000000000000000",16204 => "0000000000000000",
16205 => "0000000000000000",16206 => "0000000000000000",
16207 => "0000000000000000",16208 => "0000000000000000",
16209 => "0000000000000000",16210 => "0000000000000000",
16211 => "0000000000000000",16212 => "0000000000000000",
16213 => "0000000000000000",16214 => "0000000000000000",
16215 => "0000000000000000",16216 => "0000000000000000",
16217 => "0000000000000000",16218 => "0000000000000000",
16219 => "0000000000000000",16220 => "0000000000000000",
16221 => "0000000000000000",16222 => "0000000000000000",
16223 => "0000000000000000",16224 => "0000000000000000",
16225 => "0000000000000000",16226 => "0000000000000000",
16227 => "0000000000000000",16228 => "0000000000000000",
16229 => "0000000000000000",16230 => "0000000000000000",
16231 => "0000000000000000",16232 => "0000000000000000",
16233 => "0000000000000000",16234 => "0000000000000000",
16235 => "0000000000000000",16236 => "0000000000000000",
16237 => "0000000000000000",16238 => "0000000000000000",
16239 => "0000000000000000",16240 => "0000000000000000",
16241 => "0000000000000000",16242 => "0000000000000000",
16243 => "0000000000000000",16244 => "0000000000000000",
16245 => "0000000000000000",16246 => "0000000000000000",
16247 => "0000000000000000",16248 => "0000000000000000",
16249 => "0000000000000000",16250 => "0000000000000000",
16251 => "0000000000000000",16252 => "0000000000000000",
16253 => "0000000000000000",16254 => "0000000000000000",
16255 => "0000000000000000",16256 => "0000000000000000",
16257 => "0000000000000000",16258 => "0000000000000000",
16259 => "0000000000000000",16260 => "0000000000000000",
16261 => "0000000000000000",16262 => "0000000000000000",
16263 => "0000000000000000",16264 => "0000000000000000",
16265 => "0000000000000000",16266 => "0000000000000000",
16267 => "0000000000000000",16268 => "0000000000000000",
16269 => "0000000000000000",16270 => "0000000000000000",
16271 => "0000000000000000",16272 => "0000000000000000",
16273 => "0000000000000000",16274 => "0000000000000000",
16275 => "0000000000000000",16276 => "0000000000000000",
16277 => "0000000000000000",16278 => "0000000000000000",
16279 => "0000000000000000",16280 => "0000000000000000",
16281 => "0000000000000000",16282 => "0000000000000000",
16283 => "0000000000000000",16284 => "0000000000000000",
16285 => "0000000000000000",16286 => "0000000000000000",
16287 => "0000000000000000",16288 => "0000000000000000",
16289 => "0000000000000000",16290 => "0000000000000000",
16291 => "0000000000000000",16292 => "0000000000000000",
16293 => "0000000000000000",16294 => "0000000000000000",
16295 => "0000000000000000",16296 => "0000000000000000",
16297 => "0000000000000000",16298 => "0000000000000000",
16299 => "0000000000000000",16300 => "0000000000000000",
16301 => "0000000000000000",16302 => "0000000000000000",
16303 => "0000000000000000",16304 => "0000000000000000",
16305 => "0000000000000000",16306 => "0000000000000000",
16307 => "0000000000000000",16308 => "0000000000000000",
16309 => "0000000000000000",16310 => "0000000000000000",
16311 => "0000000000000000",16312 => "0000000000000000",
16313 => "0000000000000000",16314 => "0000000000000000",
16315 => "0000000000000000",16316 => "0000000000000000",
16317 => "0000000000000000",16318 => "0000000000000000",
16319 => "0000000000000000",16320 => "0000000000000000",
16321 => "0000000000000000",16322 => "0000000000000000",
16323 => "0000000000000000",16324 => "0000000000000000",
16325 => "0000000000000000",16326 => "0000000000000000",
16327 => "0000000000000000",16328 => "0000000000000000",
16329 => "0000000000000000",16330 => "0000000000000000",
16331 => "0000000000000000",16332 => "0000000000000000",
16333 => "0000000000000000",16334 => "0000000000000000",
16335 => "0000000000000000",16336 => "0000000000000000",
16337 => "0000000000000000",16338 => "0000000000000000",
16339 => "0000000000000000",16340 => "0000000000000000",
16341 => "0000000000000000",16342 => "0000000000000000",
16343 => "0000000000000000",16344 => "0000000000000000",
16345 => "0000000000000000",16346 => "0000000000000000",
16347 => "0000000000000000",16348 => "0000000000000000",
16349 => "0000000000000000",16350 => "0000000000000000",
16351 => "0000000000000000",16352 => "0000000000000000",
16353 => "0000000000000000",16354 => "0000000000000000",
16355 => "0000000000000000",16356 => "0000000000000000",
16357 => "0000000000000000",16358 => "0000000000000000",
16359 => "0000000000000000",16360 => "0000000000000000",
16361 => "0000000000000000",16362 => "0000000000000000",
16363 => "0000000000000000",16364 => "0000000000000000",
16365 => "0000000000000000",16366 => "0000000000000000",
16367 => "0000000000000000",16368 => "0000000000000000",
16369 => "0000000000000000",16370 => "0000000000000000",
16371 => "0000000000000000",16372 => "0000000000000000",
16373 => "0000000000000000",16374 => "0000000000000000",
16375 => "0000000000000000",16376 => "0000000000000000",
16377 => "0000000000000000",16378 => "0000000000000000",
16379 => "0000000000000000",16380 => "0000000000000000",
16381 => "0000000000000000",16382 => "0000000000000000",
16383 => "0000000000000000",16384 => "0000000000000000",
16385 => "0000000000000000",16386 => "0000000000000000",
16387 => "0000000000000000",16388 => "0000000000000000",
16389 => "0000000000000000",16390 => "0000000000000000",
16391 => "0000000000000000",16392 => "0000000000000000",
16393 => "0000000000000000",16394 => "0000000000000000",
16395 => "0000000000000000",16396 => "0000000000000000",
16397 => "0000000000000000",16398 => "0000000000000000",
16399 => "0000000000000000",16400 => "0000000000000000",
16401 => "0000000000000000",16402 => "0000000000000000",
16403 => "0000000000000000",16404 => "0000000000000000",
16405 => "0000000000000000",16406 => "0000000000000000",
16407 => "0000000000000000",16408 => "0000000000000000",
16409 => "0000000000000000",16410 => "0000000000000000",
16411 => "0000000000000000",16412 => "0000000000000000",
16413 => "0000000000000000",16414 => "0000000000000000",
16415 => "0000000000000000",16416 => "0000000000000000",
16417 => "0000000000000000",16418 => "0000000000000000",
16419 => "0000000000000000",16420 => "0000000000000000",
16421 => "0000000000000000",16422 => "0000000000000000",
16423 => "0000000000000000",16424 => "0000000000000000",
16425 => "0000000000000000",16426 => "0000000000000000",
16427 => "0000000000000000",16428 => "0000000000000000",
16429 => "0000000000000000",16430 => "0000000000000000",
16431 => "0000000000000000",16432 => "0000000000000000",
16433 => "0000000000000000",16434 => "0000000000000000",
16435 => "0000000000000000",16436 => "0000000000000000",
16437 => "0000000000000000",16438 => "0000000000000000",
16439 => "0000000000000000",16440 => "0000000000000000",
16441 => "0000000000000000",16442 => "0000000000000000",
16443 => "0000000000000000",16444 => "0000000000000000",
16445 => "0000000000000000",16446 => "0000000000000000",
16447 => "0000000000000000",16448 => "0000000000000000",
16449 => "0000000000000000",16450 => "0000000000000000",
16451 => "0000000000000000",16452 => "0000000000000000",
16453 => "0000000000000000",16454 => "0000000000000000",
16455 => "0000000000000000",16456 => "0000000000000000",
16457 => "0000000000000000",16458 => "0000000000000000",
16459 => "0000000000000000",16460 => "0000000000000000",
16461 => "0000000000000000",16462 => "0000000000000000",
16463 => "0000000000000000",16464 => "0000000000000000",
16465 => "0000000000000000",16466 => "0000000000000000",
16467 => "0000000000000000",16468 => "0000000000000000",
16469 => "0000000000000000",16470 => "0000000000000000",
16471 => "0000000000000000",16472 => "0000000000000000",
16473 => "0000000000000000",16474 => "0000000000000000",
16475 => "0000000000000000",16476 => "0000000000000000",
16477 => "0000000000000000",16478 => "0000000000000000",
16479 => "0000000000000000",16480 => "0000000000000000",
16481 => "0000000000000000",16482 => "0000000000000000",
16483 => "0000000000000000",16484 => "0000000000000000",
16485 => "0000000000000000",16486 => "0000000000000000",
16487 => "0000000000000000",16488 => "0000000000000000",
16489 => "0000000000000000",16490 => "0000000000000000",
16491 => "0000000000000000",16492 => "0000000000000000",
16493 => "0000000000000000",16494 => "0000000000000000",
16495 => "0000000000000000",16496 => "0000000000000000",
16497 => "0000000000000000",16498 => "0000000000000000",
16499 => "0000000000000000",16500 => "0000000000000000",
16501 => "0000000000000000",16502 => "0000000000000000",
16503 => "0000000000000000",16504 => "0000000000000000",
16505 => "0000000000000000",16506 => "0000000000000000",
16507 => "0000000000000000",16508 => "0000000000000000",
16509 => "0000000000000000",16510 => "0000000000000000",
16511 => "0000000000000000",16512 => "0000000000000000",
16513 => "0000000000000000",16514 => "0000000000000000",
16515 => "0000000000000000",16516 => "0000000000000000",
16517 => "0000000000000000",16518 => "0000000000000000",
16519 => "0000000000000000",16520 => "0000000000000000",
16521 => "0000000000000000",16522 => "0000000000000000",
16523 => "0000000000000000",16524 => "0000000000000000",
16525 => "0000000000000000",16526 => "0000000000000000",
16527 => "0000000000000000",16528 => "0000000000000000",
16529 => "0000000000000000",16530 => "0000000000000000",
16531 => "0000000000000000",16532 => "0000000000000000",
16533 => "0000000000000000",16534 => "0000000000000000",
16535 => "0000000000000000",16536 => "0000000000000000",
16537 => "0000000000000000",16538 => "0000000000000000",
16539 => "0000000000000000",16540 => "0000000000000000",
16541 => "0000000000000000",16542 => "0000000000000000",
16543 => "0000000000000000",16544 => "0000000000000000",
16545 => "0000000000000000",16546 => "0000000000000000",
16547 => "0000000000000000",16548 => "0000000000000000",
16549 => "0000000000000000",16550 => "0000000000000000",
16551 => "0000000000000000",16552 => "0000000000000000",
16553 => "0000000000000000",16554 => "0000000000000000",
16555 => "0000000000000000",16556 => "0000000000000000",
16557 => "0000000000000000",16558 => "0000000000000000",
16559 => "0000000000000000",16560 => "0000000000000000",
16561 => "0000000000000000",16562 => "0000000000000000",
16563 => "0000000000000000",16564 => "0000000000000000",
16565 => "0000000000000000",16566 => "0000000000000000",
16567 => "0000000000000000",16568 => "0000000000000000",
16569 => "0000000000000000",16570 => "0000000000000000",
16571 => "0000000000000000",16572 => "0000000000000000",
16573 => "0000000000000000",16574 => "0000000000000000",
16575 => "0000000000000000",16576 => "0000000000000000",
16577 => "0000000000000000",16578 => "0000000000000000",
16579 => "0000000000000000",16580 => "0000000000000000",
16581 => "0000000000000000",16582 => "0000000000000000",
16583 => "0000000000000000",16584 => "0000000000000000",
16585 => "0000000000000000",16586 => "0000000000000000",
16587 => "0000000000000000",16588 => "0000000000000000",
16589 => "0000000000000000",16590 => "0000000000000000",
16591 => "0000000000000000",16592 => "0000000000000000",
16593 => "0000000000000000",16594 => "0000000000000000",
16595 => "0000000000000000",16596 => "0000000000000000",
16597 => "0000000000000000",16598 => "0000000000000000",
16599 => "0000000000000000",16600 => "0000000000000000",
16601 => "0000000000000000",16602 => "0000000000000000",
16603 => "0000000000000000",16604 => "0000000000000000",
16605 => "0000000000000000",16606 => "0000000000000000",
16607 => "0000000000000000",16608 => "0000000000000000",
16609 => "0000000000000000",16610 => "0000000000000000",
16611 => "0000000000000000",16612 => "0000000000000000",
16613 => "0000000000000000",16614 => "0000000000000000",
16615 => "0000000000000000",16616 => "0000000000000000",
16617 => "0000000000000000",16618 => "0000000000000000",
16619 => "0000000000000000",16620 => "0000000000000000",
16621 => "0000000000000000",16622 => "0000000000000000",
16623 => "0000000000000000",16624 => "0000000000000000",
16625 => "0000000000000000",16626 => "0000000000000000",
16627 => "0000000000000000",16628 => "0000000000000000",
16629 => "0000000000000000",16630 => "0000000000000000",
16631 => "0000000000000000",16632 => "0000000000000000",
16633 => "0000000000000000",16634 => "0000000000000000",
16635 => "0000000000000000",16636 => "0000000000000000",
16637 => "0000000000000000",16638 => "0000000000000000",
16639 => "0000000000000000",16640 => "0000000000000000",
16641 => "0000000000000000",16642 => "0000000000000000",
16643 => "0000000000000000",16644 => "0000000000000000",
16645 => "0000000000000000",16646 => "0000000000000000",
16647 => "0000000000000000",16648 => "0000000000000000",
16649 => "0000000000000000",16650 => "0000000000000000",
16651 => "0000000000000000",16652 => "0000000000000000",
16653 => "0000000000000000",16654 => "0000000000000000",
16655 => "0000000000000000",16656 => "0000000000000000",
16657 => "0000000000000000",16658 => "0000000000000000",
16659 => "0000000000000000",16660 => "0000000000000000",
16661 => "0000000000000000",16662 => "0000000000000000",
16663 => "0000000000000000",16664 => "0000000000000000",
16665 => "0000000000000000",16666 => "0000000000000000",
16667 => "0000000000000000",16668 => "0000000000000000",
16669 => "0000000000000000",16670 => "0000000000000000",
16671 => "0000000000000000",16672 => "0000000000000000",
16673 => "0000000000000000",16674 => "0000000000000000",
16675 => "0000000000000000",16676 => "0000000000000000",
16677 => "0000000000000000",16678 => "0000000000000000",
16679 => "0000000000000000",16680 => "0000000000000000",
16681 => "0000000000000000",16682 => "0000000000000000",
16683 => "0000000000000000",16684 => "0000000000000000",
16685 => "0000000000000000",16686 => "0000000000000000",
16687 => "0000000000000000",16688 => "0000000000000000",
16689 => "0000000000000000",16690 => "0000000000000000",
16691 => "0000000000000000",16692 => "0000000000000000",
16693 => "0000000000000000",16694 => "0000000000000000",
16695 => "0000000000000000",16696 => "0000000000000000",
16697 => "0000000000000000",16698 => "0000000000000000",
16699 => "0000000000000000",16700 => "0000000000000000",
16701 => "0000000000000000",16702 => "0000000000000000",
16703 => "0000000000000000",16704 => "0000000000000000",
16705 => "0000000000000000",16706 => "0000000000000000",
16707 => "0000000000000000",16708 => "0000000000000000",
16709 => "0000000000000000",16710 => "0000000000000000",
16711 => "0000000000000000",16712 => "0000000000000000",
16713 => "0000000000000000",16714 => "0000000000000000",
16715 => "0000000000000000",16716 => "0000000000000000",
16717 => "0000000000000000",16718 => "0000000000000000",
16719 => "0000000000000000",16720 => "0000000000000000",
16721 => "0000000000000000",16722 => "0000000000000000",
16723 => "0000000000000000",16724 => "0000000000000000",
16725 => "0000000000000000",16726 => "0000000000000000",
16727 => "0000000000000000",16728 => "0000000000000000",
16729 => "0000000000000000",16730 => "0000000000000000",
16731 => "0000000000000000",16732 => "0000000000000000",
16733 => "0000000000000000",16734 => "0000000000000000",
16735 => "0000000000000000",16736 => "0000000000000000",
16737 => "0000000000000000",16738 => "0000000000000000",
16739 => "0000000000000000",16740 => "0000000000000000",
16741 => "0000000000000000",16742 => "0000000000000000",
16743 => "0000000000000000",16744 => "0000000000000000",
16745 => "0000000000000000",16746 => "0000000000000000",
16747 => "0000000000000000",16748 => "0000000000000000",
16749 => "0000000000000000",16750 => "0000000000000000",
16751 => "0000000000000000",16752 => "0000000000000000",
16753 => "0000000000000000",16754 => "0000000000000000",
16755 => "0000000000000000",16756 => "0000000000000000",
16757 => "0000000000000000",16758 => "0000000000000000",
16759 => "0000000000000000",16760 => "0000000000000000",
16761 => "0000000000000000",16762 => "0000000000000000",
16763 => "0000000000000000",16764 => "0000000000000000",
16765 => "0000000000000000",16766 => "0000000000000000",
16767 => "0000000000000000",16768 => "0000000000000000",
16769 => "0000000000000000",16770 => "0000000000000000",
16771 => "0000000000000000",16772 => "0000000000000000",
16773 => "0000000000000000",16774 => "0000000000000000",
16775 => "0000000000000000",16776 => "0000000000000000",
16777 => "0000000000000000",16778 => "0000000000000000",
16779 => "0000000000000000",16780 => "0000000000000000",
16781 => "0000000000000000",16782 => "0000000000000000",
16783 => "0000000000000000",16784 => "0000000000000000",
16785 => "0000000000000000",16786 => "0000000000000000",
16787 => "0000000000000000",16788 => "0000000000000000",
16789 => "0000000000000000",16790 => "0000000000000000",
16791 => "0000000000000000",16792 => "0000000000000000",
16793 => "0000000000000000",16794 => "0000000000000000",
16795 => "0000000000000000",16796 => "0000000000000000",
16797 => "0000000000000000",16798 => "0000000000000000",
16799 => "0000000000000000",16800 => "0000000000000000",
16801 => "0000000000000000",16802 => "0000000000000000",
16803 => "0000000000000000",16804 => "0000000000000000",
16805 => "0000000000000000",16806 => "0000000000000000",
16807 => "0000000000000000",16808 => "0000000000000000",
16809 => "0000000000000000",16810 => "0000000000000000",
16811 => "0000000000000000",16812 => "0000000000000000",
16813 => "0000000000000000",16814 => "0000000000000000",
16815 => "0000000000000000",16816 => "0000000000000000",
16817 => "0000000000000000",16818 => "0000000000000000",
16819 => "0000000000000000",16820 => "0000000000000000",
16821 => "0000000000000000",16822 => "0000000000000000",
16823 => "0000000000000000",16824 => "0000000000000000",
16825 => "0000000000000000",16826 => "0000000000000000",
16827 => "0000000000000000",16828 => "0000000000000000",
16829 => "0000000000000000",16830 => "0000000000000000",
16831 => "0000000000000000",16832 => "0000000000000000",
16833 => "0000000000000000",16834 => "0000000000000000",
16835 => "0000000000000000",16836 => "0000000000000000",
16837 => "0000000000000000",16838 => "0000000000000000",
16839 => "0000000000000000",16840 => "0000000000000000",
16841 => "0000000000000000",16842 => "0000000000000000",
16843 => "0000000000000000",16844 => "0000000000000000",
16845 => "0000000000000000",16846 => "0000000000000000",
16847 => "0000000000000000",16848 => "0000000000000000",
16849 => "0000000000000000",16850 => "0000000000000000",
16851 => "0000000000000000",16852 => "0000000000000000",
16853 => "0000000000000000",16854 => "0000000000000000",
16855 => "0000000000000000",16856 => "0000000000000000",
16857 => "0000000000000000",16858 => "0000000000000000",
16859 => "0000000000000000",16860 => "0000000000000000",
16861 => "0000000000000000",16862 => "0000000000000000",
16863 => "0000000000000000",16864 => "0000000000000000",
16865 => "0000000000000000",16866 => "0000000000000000",
16867 => "0000000000000000",16868 => "0000000000000000",
16869 => "0000000000000000",16870 => "0000000000000000",
16871 => "0000000000000000",16872 => "0000000000000000",
16873 => "0000000000000000",16874 => "0000000000000000",
16875 => "0000000000000000",16876 => "0000000000000000",
16877 => "0000000000000000",16878 => "0000000000000000",
16879 => "0000000000000000",16880 => "0000000000000000",
16881 => "0000000000000000",16882 => "0000000000000000",
16883 => "0000000000000000",16884 => "0000000000000000",
16885 => "0000000000000000",16886 => "0000000000000000",
16887 => "0000000000000000",16888 => "0000000000000000",
16889 => "0000000000000000",16890 => "0000000000000000",
16891 => "0000000000000000",16892 => "0000000000000000",
16893 => "0000000000000000",16894 => "0000000000000000",
16895 => "0000000000000000",16896 => "0000000000000000",
16897 => "0000000000000000",16898 => "0000000000000000",
16899 => "0000000000000000",16900 => "0000000000000000",
16901 => "0000000000000000",16902 => "0000000000000000",
16903 => "0000000000000000",16904 => "0000000000000000",
16905 => "0000000000000000",16906 => "0000000000000000",
16907 => "0000000000000000",16908 => "0000000000000000",
16909 => "0000000000000000",16910 => "0000000000000000",
16911 => "0000000000000000",16912 => "0000000000000000",
16913 => "0000000000000000",16914 => "0000000000000000",
16915 => "0000000000000000",16916 => "0000000000000000",
16917 => "0000000000000000",16918 => "0000000000000000",
16919 => "0000000000000000",16920 => "0000000000000000",
16921 => "0000000000000000",16922 => "0000000000000000",
16923 => "0000000000000000",16924 => "0000000000000000",
16925 => "0000000000000000",16926 => "0000000000000000",
16927 => "0000000000000000",16928 => "0000000000000000",
16929 => "0000000000000000",16930 => "0000000000000000",
16931 => "0000000000000000",16932 => "0000000000000000",
16933 => "0000000000000000",16934 => "0000000000000000",
16935 => "0000000000000000",16936 => "0000000000000000",
16937 => "0000000000000000",16938 => "0000000000000000",
16939 => "0000000000000000",16940 => "0000000000000000",
16941 => "0000000000000000",16942 => "0000000000000000",
16943 => "0000000000000000",16944 => "0000000000000000",
16945 => "0000000000000000",16946 => "0000000000000000",
16947 => "0000000000000000",16948 => "0000000000000000",
16949 => "0000000000000000",16950 => "0000000000000000",
16951 => "0000000000000000",16952 => "0000000000000000",
16953 => "0000000000000000",16954 => "0000000000000000",
16955 => "0000000000000000",16956 => "0000000000000000",
16957 => "0000000000000000",16958 => "0000000000000000",
16959 => "0000000000000000",16960 => "0000000000000000",
16961 => "0000000000000000",16962 => "0000000000000000",
16963 => "0000000000000000",16964 => "0000000000000000",
16965 => "0000000000000000",16966 => "0000000000000000",
16967 => "0000000000000000",16968 => "0000000000000000",
16969 => "0000000000000000",16970 => "0000000000000000",
16971 => "0000000000000000",16972 => "0000000000000000",
16973 => "0000000000000000",16974 => "0000000000000000",
16975 => "0000000000000000",16976 => "0000000000000000",
16977 => "0000000000000000",16978 => "0000000000000000",
16979 => "0000000000000000",16980 => "0000000000000000",
16981 => "0000000000000000",16982 => "0000000000000000",
16983 => "0000000000000000",16984 => "0000000000000000",
16985 => "0000000000000000",16986 => "0000000000000000",
16987 => "0000000000000000",16988 => "0000000000000000",
16989 => "0000000000000000",16990 => "0000000000000000",
16991 => "0000000000000000",16992 => "0000000000000000",
16993 => "0000000000000000",16994 => "0000000000000000",
16995 => "0000000000000000",16996 => "0000000000000000",
16997 => "0000000000000000",16998 => "0000000000000000",
16999 => "0000000000000000",17000 => "0000000000000000",
17001 => "0000000000000000",17002 => "0000000000000000",
17003 => "0000000000000000",17004 => "0000000000000000",
17005 => "0000000000000000",17006 => "0000000000000000",
17007 => "0000000000000000",17008 => "0000000000000000",
17009 => "0000000000000000",17010 => "0000000000000000",
17011 => "0000000000000000",17012 => "0000000000000000",
17013 => "0000000000000000",17014 => "0000000000000000",
17015 => "0000000000000000",17016 => "0000000000000000",
17017 => "0000000000000000",17018 => "0000000000000000",
17019 => "0000000000000000",17020 => "0000000000000000",
17021 => "0000000000000000",17022 => "0000000000000000",
17023 => "0000000000000000",17024 => "0000000000000000",
17025 => "0000000000000000",17026 => "0000000000000000",
17027 => "0000000000000000",17028 => "0000000000000000",
17029 => "0000000000000000",17030 => "0000000000000000",
17031 => "0000000000000000",17032 => "0000000000000000",
17033 => "0000000000000000",17034 => "0000000000000000",
17035 => "0000000000000000",17036 => "0000000000000000",
17037 => "0000000000000000",17038 => "0000000000000000",
17039 => "0000000000000000",17040 => "0000000000000000",
17041 => "0000000000000000",17042 => "0000000000000000",
17043 => "0000000000000000",17044 => "0000000000000000",
17045 => "0000000000000000",17046 => "0000000000000000",
17047 => "0000000000000000",17048 => "0000000000000000",
17049 => "0000000000000000",17050 => "0000000000000000",
17051 => "0000000000000000",17052 => "0000000000000000",
17053 => "0000000000000000",17054 => "0000000000000000",
17055 => "0000000000000000",17056 => "0000000000000000",
17057 => "0000000000000000",17058 => "0000000000000000",
17059 => "0000000000000000",17060 => "0000000000000000",
17061 => "0000000000000000",17062 => "0000000000000000",
17063 => "0000000000000000",17064 => "0000000000000000",
17065 => "0000000000000000",17066 => "0000000000000000",
17067 => "0000000000000000",17068 => "0000000000000000",
17069 => "0000000000000000",17070 => "0000000000000000",
17071 => "0000000000000000",17072 => "0000000000000000",
17073 => "0000000000000000",17074 => "0000000000000000",
17075 => "0000000000000000",17076 => "0000000000000000",
17077 => "0000000000000000",17078 => "0000000000000000",
17079 => "0000000000000000",17080 => "0000000000000000",
17081 => "0000000000000000",17082 => "0000000000000000",
17083 => "0000000000000000",17084 => "0000000000000000",
17085 => "0000000000000000",17086 => "0000000000000000",
17087 => "0000000000000000",17088 => "0000000000000000",
17089 => "0000000000000000",17090 => "0000000000000000",
17091 => "0000000000000000",17092 => "0000000000000000",
17093 => "0000000000000000",17094 => "0000000000000000",
17095 => "0000000000000000",17096 => "0000000000000000",
17097 => "0000000000000000",17098 => "0000000000000000",
17099 => "0000000000000000",17100 => "0000000000000000",
17101 => "0000000000000000",17102 => "0000000000000000",
17103 => "0000000000000000",17104 => "0000000000000000",
17105 => "0000000000000000",17106 => "0000000000000000",
17107 => "0000000000000000",17108 => "0000000000000000",
17109 => "0000000000000000",17110 => "0000000000000000",
17111 => "0000000000000000",17112 => "0000000000000000",
17113 => "0000000000000000",17114 => "0000000000000000",
17115 => "0000000000000000",17116 => "0000000000000000",
17117 => "0000000000000000",17118 => "0000000000000000",
17119 => "0000000000000000",17120 => "0000000000000000",
17121 => "0000000000000000",17122 => "0000000000000000",
17123 => "0000000000000000",17124 => "0000000000000000",
17125 => "0000000000000000",17126 => "0000000000000000",
17127 => "0000000000000000",17128 => "0000000000000000",
17129 => "0000000000000000",17130 => "0000000000000000",
17131 => "0000000000000000",17132 => "0000000000000000",
17133 => "0000000000000000",17134 => "0000000000000000",
17135 => "0000000000000000",17136 => "0000000000000000",
17137 => "0000000000000000",17138 => "0000000000000000",
17139 => "0000000000000000",17140 => "0000000000000000",
17141 => "0000000000000000",17142 => "0000000000000000",
17143 => "0000000000000000",17144 => "0000000000000000",
17145 => "0000000000000000",17146 => "0000000000000000",
17147 => "0000000000000000",17148 => "0000000000000000",
17149 => "0000000000000000",17150 => "0000000000000000",
17151 => "0000000000000000",17152 => "0000000000000000",
17153 => "0000000000000000",17154 => "0000000000000000",
17155 => "0000000000000000",17156 => "0000000000000000",
17157 => "0000000000000000",17158 => "0000000000000000",
17159 => "0000000000000000",17160 => "0000000000000000",
17161 => "0000000000000000",17162 => "0000000000000000",
17163 => "0000000000000000",17164 => "0000000000000000",
17165 => "0000000000000000",17166 => "0000000000000000",
17167 => "0000000000000000",17168 => "0000000000000000",
17169 => "0000000000000000",17170 => "0000000000000000",
17171 => "0000000000000000",17172 => "0000000000000000",
17173 => "0000000000000000",17174 => "0000000000000000",
17175 => "0000000000000000",17176 => "0000000000000000",
17177 => "0000000000000000",17178 => "0000000000000000",
17179 => "0000000000000000",17180 => "0000000000000000",
17181 => "0000000000000000",17182 => "0000000000000000",
17183 => "0000000000000000",17184 => "0000000000000000",
17185 => "0000000000000000",17186 => "0000000000000000",
17187 => "0000000000000000",17188 => "0000000000000000",
17189 => "0000000000000000",17190 => "0000000000000000",
17191 => "0000000000000000",17192 => "0000000000000000",
17193 => "0000000000000000",17194 => "0000000000000000",
17195 => "0000000000000000",17196 => "0000000000000000",
17197 => "0000000000000000",17198 => "0000000000000000",
17199 => "0000000000000000",17200 => "0000000000000000",
17201 => "0000000000000000",17202 => "0000000000000000",
17203 => "0000000000000000",17204 => "0000000000000000",
17205 => "0000000000000000",17206 => "0000000000000000",
17207 => "0000000000000000",17208 => "0000000000000000",
17209 => "0000000000000000",17210 => "0000000000000000",
17211 => "0000000000000000",17212 => "0000000000000000",
17213 => "0000000000000000",17214 => "0000000000000000",
17215 => "0000000000000000",17216 => "0000000000000000",
17217 => "0000000000000000",17218 => "0000000000000000",
17219 => "0000000000000000",17220 => "0000000000000000",
17221 => "0000000000000000",17222 => "0000000000000000",
17223 => "0000000000000000",17224 => "0000000000000000",
17225 => "0000000000000000",17226 => "0000000000000000",
17227 => "0000000000000000",17228 => "0000000000000000",
17229 => "0000000000000000",17230 => "0000000000000000",
17231 => "0000000000000000",17232 => "0000000000000000",
17233 => "0000000000000000",17234 => "0000000000000000",
17235 => "0000000000000000",17236 => "0000000000000000",
17237 => "0000000000000000",17238 => "0000000000000000",
17239 => "0000000000000000",17240 => "0000000000000000",
17241 => "0000000000000000",17242 => "0000000000000000",
17243 => "0000000000000000",17244 => "0000000000000000",
17245 => "0000000000000000",17246 => "0000000000000000",
17247 => "0000000000000000",17248 => "0000000000000000",
17249 => "0000000000000000",17250 => "0000000000000000",
17251 => "0000000000000000",17252 => "0000000000000000",
17253 => "0000000000000000",17254 => "0000000000000000",
17255 => "0000000000000000",17256 => "0000000000000000",
17257 => "0000000000000000",17258 => "0000000000000000",
17259 => "0000000000000000",17260 => "0000000000000000",
17261 => "0000000000000000",17262 => "0000000000000000",
17263 => "0000000000000000",17264 => "0000000000000000",
17265 => "0000000000000000",17266 => "0000000000000000",
17267 => "0000000000000000",17268 => "0000000000000000",
17269 => "0000000000000000",17270 => "0000000000000000",
17271 => "0000000000000000",17272 => "0000000000000000",
17273 => "0000000000000000",17274 => "0000000000000000",
17275 => "0000000000000000",17276 => "0000000000000000",
17277 => "0000000000000000",17278 => "0000000000000000",
17279 => "0000000000000000",17280 => "0000000000000000",
17281 => "0000000000000000",17282 => "0000000000000000",
17283 => "0000000000000000",17284 => "0000000000000000",
17285 => "0000000000000000",17286 => "0000000000000000",
17287 => "0000000000000000",17288 => "0000000000000000",
17289 => "0000000000000000",17290 => "0000000000000000",
17291 => "0000000000000000",17292 => "0000000000000000",
17293 => "0000000000000000",17294 => "0000000000000000",
17295 => "0000000000000000",17296 => "0000000000000000",
17297 => "0000000000000000",17298 => "0000000000000000",
17299 => "0000000000000000",17300 => "0000000000000000",
17301 => "0000000000000000",17302 => "0000000000000000",
17303 => "0000000000000000",17304 => "0000000000000000",
17305 => "0000000000000000",17306 => "0000000000000000",
17307 => "0000000000000000",17308 => "0000000000000000",
17309 => "0000000000000000",17310 => "0000000000000000",
17311 => "0000000000000000",17312 => "0000000000000000",
17313 => "0000000000000000",17314 => "0000000000000000",
17315 => "0000000000000000",17316 => "0000000000000000",
17317 => "0000000000000000",17318 => "0000000000000000",
17319 => "0000000000000000",17320 => "0000000000000000",
17321 => "0000000000000000",17322 => "0000000000000000",
17323 => "0000000000000000",17324 => "0000000000000000",
17325 => "0000000000000000",17326 => "0000000000000000",
17327 => "0000000000000000",17328 => "0000000000000000",
17329 => "0000000000000000",17330 => "0000000000000000",
17331 => "0000000000000000",17332 => "0000000000000000",
17333 => "0000000000000000",17334 => "0000000000000000",
17335 => "0000000000000000",17336 => "0000000000000000",
17337 => "0000000000000000",17338 => "0000000000000000",
17339 => "0000000000000000",17340 => "0000000000000000",
17341 => "0000000000000000",17342 => "0000000000000000",
17343 => "0000000000000000",17344 => "0000000000000000",
17345 => "0000000000000000",17346 => "0000000000000000",
17347 => "0000000000000000",17348 => "0000000000000000",
17349 => "0000000000000000",17350 => "0000000000000000",
17351 => "0000000000000000",17352 => "0000000000000000",
17353 => "0000000000000000",17354 => "0000000000000000",
17355 => "0000000000000000",17356 => "0000000000000000",
17357 => "0000000000000000",17358 => "0000000000000000",
17359 => "0000000000000000",17360 => "0000000000000000",
17361 => "0000000000000000",17362 => "0000000000000000",
17363 => "0000000000000000",17364 => "0000000000000000",
17365 => "0000000000000000",17366 => "0000000000000000",
17367 => "0000000000000000",17368 => "0000000000000000",
17369 => "0000000000000000",17370 => "0000000000000000",
17371 => "0000000000000000",17372 => "0000000000000000",
17373 => "0000000000000000",17374 => "0000000000000000",
17375 => "0000000000000000",17376 => "0000000000000000",
17377 => "0000000000000000",17378 => "0000000000000000",
17379 => "0000000000000000",17380 => "0000000000000000",
17381 => "0000000000000000",17382 => "0000000000000000",
17383 => "0000000000000000",17384 => "0000000000000000",
17385 => "0000000000000000",17386 => "0000000000000000",
17387 => "0000000000000000",17388 => "0000000000000000",
17389 => "0000000000000000",17390 => "0000000000000000",
17391 => "0000000000000000",17392 => "0000000000000000",
17393 => "0000000000000000",17394 => "0000000000000000",
17395 => "0000000000000000",17396 => "0000000000000000",
17397 => "0000000000000000",17398 => "0000000000000000",
17399 => "0000000000000000",17400 => "0000000000000000",
17401 => "0000000000000000",17402 => "0000000000000000",
17403 => "0000000000000000",17404 => "0000000000000000",
17405 => "0000000000000000",17406 => "0000000000000000",
17407 => "0000000000000000",17408 => "0000000000000000",
17409 => "0000000000000000",17410 => "0000000000000000",
17411 => "0000000000000000",17412 => "0000000000000000",
17413 => "0000000000000000",17414 => "0000000000000000",
17415 => "0000000000000000",17416 => "0000000000000000",
17417 => "0000000000000000",17418 => "0000000000000000",
17419 => "0000000000000000",17420 => "0000000000000000",
17421 => "0000000000000000",17422 => "0000000000000000",
17423 => "0000000000000000",17424 => "0000000000000000",
17425 => "0000000000000000",17426 => "0000000000000000",
17427 => "0000000000000000",17428 => "0000000000000000",
17429 => "0000000000000000",17430 => "0000000000000000",
17431 => "0000000000000000",17432 => "0000000000000000",
17433 => "0000000000000000",17434 => "0000000000000000",
17435 => "0000000000000000",17436 => "0000000000000000",
17437 => "0000000000000000",17438 => "0000000000000000",
17439 => "0000000000000000",17440 => "0000000000000000",
17441 => "0000000000000000",17442 => "0000000000000000",
17443 => "0000000000000000",17444 => "0000000000000000",
17445 => "0000000000000000",17446 => "0000000000000000",
17447 => "0000000000000000",17448 => "0000000000000000",
17449 => "0000000000000000",17450 => "0000000000000000",
17451 => "0000000000000000",17452 => "0000000000000000",
17453 => "0000000000000000",17454 => "0000000000000000",
17455 => "0000000000000000",17456 => "0000000000000000",
17457 => "0000000000000000",17458 => "0000000000000000",
17459 => "0000000000000000",17460 => "0000000000000000",
17461 => "0000000000000000",17462 => "0000000000000000",
17463 => "0000000000000000",17464 => "0000000000000000",
17465 => "0000000000000000",17466 => "0000000000000000",
17467 => "0000000000000000",17468 => "0000000000000000",
17469 => "0000000000000000",17470 => "0000000000000000",
17471 => "0000000000000000",17472 => "0000000000000000",
17473 => "0000000000000000",17474 => "0000000000000000",
17475 => "0000000000000000",17476 => "0000000000000000",
17477 => "0000000000000000",17478 => "0000000000000000",
17479 => "0000000000000000",17480 => "0000000000000000",
17481 => "0000000000000000",17482 => "0000000000000000",
17483 => "0000000000000000",17484 => "0000000000000000",
17485 => "0000000000000000",17486 => "0000000000000000",
17487 => "0000000000000000",17488 => "0000000000000000",
17489 => "0000000000000000",17490 => "0000000000000000",
17491 => "0000000000000000",17492 => "0000000000000000",
17493 => "0000000000000000",17494 => "0000000000000000",
17495 => "0000000000000000",17496 => "0000000000000000",
17497 => "0000000000000000",17498 => "0000000000000000",
17499 => "0000000000000000",17500 => "0000000000000000",
17501 => "0000000000000000",17502 => "0000000000000000",
17503 => "0000000000000000",17504 => "0000000000000000",
17505 => "0000000000000000",17506 => "0000000000000000",
17507 => "0000000000000000",17508 => "0000000000000000",
17509 => "0000000000000000",17510 => "0000000000000000",
17511 => "0000000000000000",17512 => "0000000000000000",
17513 => "0000000000000000",17514 => "0000000000000000",
17515 => "0000000000000000",17516 => "0000000000000000",
17517 => "0000000000000000",17518 => "0000000000000000",
17519 => "0000000000000000",17520 => "0000000000000000",
17521 => "0000000000000000",17522 => "0000000000000000",
17523 => "0000000000000000",17524 => "0000000000000000",
17525 => "0000000000000000",17526 => "0000000000000000",
17527 => "0000000000000000",17528 => "0000000000000000",
17529 => "0000000000000000",17530 => "0000000000000000",
17531 => "0000000000000000",17532 => "0000000000000000",
17533 => "0000000000000000",17534 => "0000000000000000",
17535 => "0000000000000000",17536 => "0000000000000000",
17537 => "0000000000000000",17538 => "0000000000000000",
17539 => "0000000000000000",17540 => "0000000000000000",
17541 => "0000000000000000",17542 => "0000000000000000",
17543 => "0000000000000000",17544 => "0000000000000000",
17545 => "0000000000000000",17546 => "0000000000000000",
17547 => "0000000000000000",17548 => "0000000000000000",
17549 => "0000000000000000",17550 => "0000000000000000",
17551 => "0000000000000000",17552 => "0000000000000000",
17553 => "0000000000000000",17554 => "0000000000000000",
17555 => "0000000000000000",17556 => "0000000000000000",
17557 => "0000000000000000",17558 => "0000000000000000",
17559 => "0000000000000000",17560 => "0000000000000000",
17561 => "0000000000000000",17562 => "0000000000000000",
17563 => "0000000000000000",17564 => "0000000000000000",
17565 => "0000000000000000",17566 => "0000000000000000",
17567 => "0000000000000000",17568 => "0000000000000000",
17569 => "0000000000000000",17570 => "0000000000000000",
17571 => "0000000000000000",17572 => "0000000000000000",
17573 => "0000000000000000",17574 => "0000000000000000",
17575 => "0000000000000000",17576 => "0000000000000000",
17577 => "0000000000000000",17578 => "0000000000000000",
17579 => "0000000000000000",17580 => "0000000000000000",
17581 => "0000000000000000",17582 => "0000000000000000",
17583 => "0000000000000000",17584 => "0000000000000000",
17585 => "0000000000000000",17586 => "0000000000000000",
17587 => "0000000000000000",17588 => "0000000000000000",
17589 => "0000000000000000",17590 => "0000000000000000",
17591 => "0000000000000000",17592 => "0000000000000000",
17593 => "0000000000000000",17594 => "0000000000000000",
17595 => "0000000000000000",17596 => "0000000000000000",
17597 => "0000000000000000",17598 => "0000000000000000",
17599 => "0000000000000000",17600 => "0000000000000000",
17601 => "0000000000000000",17602 => "0000000000000000",
17603 => "0000000000000000",17604 => "0000000000000000",
17605 => "0000000000000000",17606 => "0000000000000000",
17607 => "0000000000000000",17608 => "0000000000000000",
17609 => "0000000000000000",17610 => "0000000000000000",
17611 => "0000000000000000",17612 => "0000000000000000",
17613 => "0000000000000000",17614 => "0000000000000000",
17615 => "0000000000000000",17616 => "0000000000000000",
17617 => "0000000000000000",17618 => "0000000000000000",
17619 => "0000000000000000",17620 => "0000000000000000",
17621 => "0000000000000000",17622 => "0000000000000000",
17623 => "0000000000000000",17624 => "0000000000000000",
17625 => "0000000000000000",17626 => "0000000000000000",
17627 => "0000000000000000",17628 => "0000000000000000",
17629 => "0000000000000000",17630 => "0000000000000000",
17631 => "0000000000000000",17632 => "0000000000000000",
17633 => "0000000000000000",17634 => "0000000000000000",
17635 => "0000000000000000",17636 => "0000000000000000",
17637 => "0000000000000000",17638 => "0000000000000000",
17639 => "0000000000000000",17640 => "0000000000000000",
17641 => "0000000000000000",17642 => "0000000000000000",
17643 => "0000000000000000",17644 => "0000000000000000",
17645 => "0000000000000000",17646 => "0000000000000000",
17647 => "0000000000000000",17648 => "0000000000000000",
17649 => "0000000000000000",17650 => "0000000000000000",
17651 => "0000000000000000",17652 => "0000000000000000",
17653 => "0000000000000000",17654 => "0000000000000000",
17655 => "0000000000000000",17656 => "0000000000000000",
17657 => "0000000000000000",17658 => "0000000000000000",
17659 => "0000000000000000",17660 => "0000000000000000",
17661 => "0000000000000000",17662 => "0000000000000000",
17663 => "0000000000000000",17664 => "0000000000000000",
17665 => "0000000000000000",17666 => "0000000000000000",
17667 => "0000000000000000",17668 => "0000000000000000",
17669 => "0000000000000000",17670 => "0000000000000000",
17671 => "0000000000000000",17672 => "0000000000000000",
17673 => "0000000000000000",17674 => "0000000000000000",
17675 => "0000000000000000",17676 => "0000000000000000",
17677 => "0000000000000000",17678 => "0000000000000000",
17679 => "0000000000000000",17680 => "0000000000000000",
17681 => "0000000000000000",17682 => "0000000000000000",
17683 => "0000000000000000",17684 => "0000000000000000",
17685 => "0000000000000000",17686 => "0000000000000000",
17687 => "0000000000000000",17688 => "0000000000000000",
17689 => "0000000000000000",17690 => "0000000000000000",
17691 => "0000000000000000",17692 => "0000000000000000",
17693 => "0000000000000000",17694 => "0000000000000000",
17695 => "0000000000000000",17696 => "0000000000000000",
17697 => "0000000000000000",17698 => "0000000000000000",
17699 => "0000000000000000",17700 => "0000000000000000",
17701 => "0000000000000000",17702 => "0000000000000000",
17703 => "0000000000000000",17704 => "0000000000000000",
17705 => "0000000000000000",17706 => "0000000000000000",
17707 => "0000000000000000",17708 => "0000000000000000",
17709 => "0000000000000000",17710 => "0000000000000000",
17711 => "0000000000000000",17712 => "0000000000000000",
17713 => "0000000000000000",17714 => "0000000000000000",
17715 => "0000000000000000",17716 => "0000000000000000",
17717 => "0000000000000000",17718 => "0000000000000000",
17719 => "0000000000000000",17720 => "0000000000000000",
17721 => "0000000000000000",17722 => "0000000000000000",
17723 => "0000000000000000",17724 => "0000000000000000",
17725 => "0000000000000000",17726 => "0000000000000000",
17727 => "0000000000000000",17728 => "0000000000000000",
17729 => "0000000000000000",17730 => "0000000000000000",
17731 => "0000000000000000",17732 => "0000000000000000",
17733 => "0000000000000000",17734 => "0000000000000000",
17735 => "0000000000000000",17736 => "0000000000000000",
17737 => "0000000000000000",17738 => "0000000000000000",
17739 => "0000000000000000",17740 => "0000000000000000",
17741 => "0000000000000000",17742 => "0000000000000000",
17743 => "0000000000000000",17744 => "0000000000000000",
17745 => "0000000000000000",17746 => "0000000000000000",
17747 => "0000000000000000",17748 => "0000000000000000",
17749 => "0000000000000000",17750 => "0000000000000000",
17751 => "0000000000000000",17752 => "0000000000000000",
17753 => "0000000000000000",17754 => "0000000000000000",
17755 => "0000000000000000",17756 => "0000000000000000",
17757 => "0000000000000000",17758 => "0000000000000000",
17759 => "0000000000000000",17760 => "0000000000000000",
17761 => "0000000000000000",17762 => "0000000000000000",
17763 => "0000000000000000",17764 => "0000000000000000",
17765 => "0000000000000000",17766 => "0000000000000000",
17767 => "0000000000000000",17768 => "0000000000000000",
17769 => "0000000000000000",17770 => "0000000000000000",
17771 => "0000000000000000",17772 => "0000000000000000",
17773 => "0000000000000000",17774 => "0000000000000000",
17775 => "0000000000000000",17776 => "0000000000000000",
17777 => "0000000000000000",17778 => "0000000000000000",
17779 => "0000000000000000",17780 => "0000000000000000",
17781 => "0000000000000000",17782 => "0000000000000000",
17783 => "0000000000000000",17784 => "0000000000000000",
17785 => "0000000000000000",17786 => "0000000000000000",
17787 => "0000000000000000",17788 => "0000000000000000",
17789 => "0000000000000000",17790 => "0000000000000000",
17791 => "0000000000000000",17792 => "0000000000000000",
17793 => "0000000000000000",17794 => "0000000000000000",
17795 => "0000000000000000",17796 => "0000000000000000",
17797 => "0000000000000000",17798 => "0000000000000000",
17799 => "0000000000000000",17800 => "0000000000000000",
17801 => "0000000000000000",17802 => "0000000000000000",
17803 => "0000000000000000",17804 => "0000000000000000",
17805 => "0000000000000000",17806 => "0000000000000000",
17807 => "0000000000000000",17808 => "0000000000000000",
17809 => "0000000000000000",17810 => "0000000000000000",
17811 => "0000000000000000",17812 => "0000000000000000",
17813 => "0000000000000000",17814 => "0000000000000000",
17815 => "0000000000000000",17816 => "0000000000000000",
17817 => "0000000000000000",17818 => "0000000000000000",
17819 => "0000000000000000",17820 => "0000000000000000",
17821 => "0000000000000000",17822 => "0000000000000000",
17823 => "0000000000000000",17824 => "0000000000000000",
17825 => "0000000000000000",17826 => "0000000000000000",
17827 => "0000000000000000",17828 => "0000000000000000",
17829 => "0000000000000000",17830 => "0000000000000000",
17831 => "0000000000000000",17832 => "0000000000000000",
17833 => "0000000000000000",17834 => "0000000000000000",
17835 => "0000000000000000",17836 => "0000000000000000",
17837 => "0000000000000000",17838 => "0000000000000000",
17839 => "0000000000000000",17840 => "0000000000000000",
17841 => "0000000000000000",17842 => "0000000000000000",
17843 => "0000000000000000",17844 => "0000000000000000",
17845 => "0000000000000000",17846 => "0000000000000000",
17847 => "0000000000000000",17848 => "0000000000000000",
17849 => "0000000000000000",17850 => "0000000000000000",
17851 => "0000000000000000",17852 => "0000000000000000",
17853 => "0000000000000000",17854 => "0000000000000000",
17855 => "0000000000000000",17856 => "0000000000000000",
17857 => "0000000000000000",17858 => "0000000000000000",
17859 => "0000000000000000",17860 => "0000000000000000",
17861 => "0000000000000000",17862 => "0000000000000000",
17863 => "0000000000000000",17864 => "0000000000000000",
17865 => "0000000000000000",17866 => "0000000000000000",
17867 => "0000000000000000",17868 => "0000000000000000",
17869 => "0000000000000000",17870 => "0000000000000000",
17871 => "0000000000000000",17872 => "0000000000000000",
17873 => "0000000000000000",17874 => "0000000000000000",
17875 => "0000000000000000",17876 => "0000000000000000",
17877 => "0000000000000000",17878 => "0000000000000000",
17879 => "0000000000000000",17880 => "0000000000000000",
17881 => "0000000000000000",17882 => "0000000000000000",
17883 => "0000000000000000",17884 => "0000000000000000",
17885 => "0000000000000000",17886 => "0000000000000000",
17887 => "0000000000000000",17888 => "0000000000000000",
17889 => "0000000000000000",17890 => "0000000000000000",
17891 => "0000000000000000",17892 => "0000000000000000",
17893 => "0000000000000000",17894 => "0000000000000000",
17895 => "0000000000000000",17896 => "0000000000000000",
17897 => "0000000000000000",17898 => "0000000000000000",
17899 => "0000000000000000",17900 => "0000000000000000",
17901 => "0000000000000000",17902 => "0000000000000000",
17903 => "0000000000000000",17904 => "0000000000000000",
17905 => "0000000000000000",17906 => "0000000000000000",
17907 => "0000000000000000",17908 => "0000000000000000",
17909 => "0000000000000000",17910 => "0000000000000000",
17911 => "0000000000000000",17912 => "0000000000000000",
17913 => "0000000000000000",17914 => "0000000000000000",
17915 => "0000000000000000",17916 => "0000000000000000",
17917 => "0000000000000000",17918 => "0000000000000000",
17919 => "0000000000000000",17920 => "0000000000000000",
17921 => "0000000000000000",17922 => "0000000000000000",
17923 => "0000000000000000",17924 => "0000000000000000",
17925 => "0000000000000000",17926 => "0000000000000000",
17927 => "0000000000000000",17928 => "0000000000000000",
17929 => "0000000000000000",17930 => "0000000000000000",
17931 => "0000000000000000",17932 => "0000000000000000",
17933 => "0000000000000000",17934 => "0000000000000000",
17935 => "0000000000000000",17936 => "0000000000000000",
17937 => "0000000000000000",17938 => "0000000000000000",
17939 => "0000000000000000",17940 => "0000000000000000",
17941 => "0000000000000000",17942 => "0000000000000000",
17943 => "0000000000000000",17944 => "0000000000000000",
17945 => "0000000000000000",17946 => "0000000000000000",
17947 => "0000000000000000",17948 => "0000000000000000",
17949 => "0000000000000000",17950 => "0000000000000000",
17951 => "0000000000000000",17952 => "0000000000000000",
17953 => "0000000000000000",17954 => "0000000000000000",
17955 => "0000000000000000",17956 => "0000000000000000",
17957 => "0000000000000000",17958 => "0000000000000000",
17959 => "0000000000000000",17960 => "0000000000000000",
17961 => "0000000000000000",17962 => "0000000000000000",
17963 => "0000000000000000",17964 => "0000000000000000",
17965 => "0000000000000000",17966 => "0000000000000000",
17967 => "0000000000000000",17968 => "0000000000000000",
17969 => "0000000000000000",17970 => "0000000000000000",
17971 => "0000000000000000",17972 => "0000000000000000",
17973 => "0000000000000000",17974 => "0000000000000000",
17975 => "0000000000000000",17976 => "0000000000000000",
17977 => "0000000000000000",17978 => "0000000000000000",
17979 => "0000000000000000",17980 => "0000000000000000",
17981 => "0000000000000000",17982 => "0000000000000000",
17983 => "0000000000000000",17984 => "0000000000000000",
17985 => "0000000000000000",17986 => "0000000000000000",
17987 => "0000000000000000",17988 => "0000000000000000",
17989 => "0000000000000000",17990 => "0000000000000000",
17991 => "0000000000000000",17992 => "0000000000000000",
17993 => "0000000000000000",17994 => "0000000000000000",
17995 => "0000000000000000",17996 => "0000000000000000",
17997 => "0000000000000000",17998 => "0000000000000000",
17999 => "0000000000000000",18000 => "0000000000000000",
18001 => "0000000000000000",18002 => "0000000000000000",
18003 => "0000000000000000",18004 => "0000000000000000",
18005 => "0000000000000000",18006 => "0000000000000000",
18007 => "0000000000000000",18008 => "0000000000000000",
18009 => "0000000000000000",18010 => "0000000000000000",
18011 => "0000000000000000",18012 => "0000000000000000",
18013 => "0000000000000000",18014 => "0000000000000000",
18015 => "0000000000000000",18016 => "0000000000000000",
18017 => "0000000000000000",18018 => "0000000000000000",
18019 => "0000000000000000",18020 => "0000000000000000",
18021 => "0000000000000000",18022 => "0000000000000000",
18023 => "0000000000000000",18024 => "0000000000000000",
18025 => "0000000000000000",18026 => "0000000000000000",
18027 => "0000000000000000",18028 => "0000000000000000",
18029 => "0000000000000000",18030 => "0000000000000000",
18031 => "0000000000000000",18032 => "0000000000000000",
18033 => "0000000000000000",18034 => "0000000000000000",
18035 => "0000000000000000",18036 => "0000000000000000",
18037 => "0000000000000000",18038 => "0000000000000000",
18039 => "0000000000000000",18040 => "0000000000000000",
18041 => "0000000000000000",18042 => "0000000000000000",
18043 => "0000000000000000",18044 => "0000000000000000",
18045 => "0000000000000000",18046 => "0000000000000000",
18047 => "0000000000000000",18048 => "0000000000000000",
18049 => "0000000000000000",18050 => "0000000000000000",
18051 => "0000000000000000",18052 => "0000000000000000",
18053 => "0000000000000000",18054 => "0000000000000000",
18055 => "0000000000000000",18056 => "0000000000000000",
18057 => "0000000000000000",18058 => "0000000000000000",
18059 => "0000000000000000",18060 => "0000000000000000",
18061 => "0000000000000000",18062 => "0000000000000000",
18063 => "0000000000000000",18064 => "0000000000000000",
18065 => "0000000000000000",18066 => "0000000000000000",
18067 => "0000000000000000",18068 => "0000000000000000",
18069 => "0000000000000000",18070 => "0000000000000000",
18071 => "0000000000000000",18072 => "0000000000000000",
18073 => "0000000000000000",18074 => "0000000000000000",
18075 => "0000000000000000",18076 => "0000000000000000",
18077 => "0000000000000000",18078 => "0000000000000000",
18079 => "0000000000000000",18080 => "0000000000000000",
18081 => "0000000000000000",18082 => "0000000000000000",
18083 => "0000000000000000",18084 => "0000000000000000",
18085 => "0000000000000000",18086 => "0000000000000000",
18087 => "0000000000000000",18088 => "0000000000000000",
18089 => "0000000000000000",18090 => "0000000000000000",
18091 => "0000000000000000",18092 => "0000000000000000",
18093 => "0000000000000000",18094 => "0000000000000000",
18095 => "0000000000000000",18096 => "0000000000000000",
18097 => "0000000000000000",18098 => "0000000000000000",
18099 => "0000000000000000",18100 => "0000000000000000",
18101 => "0000000000000000",18102 => "0000000000000000",
18103 => "0000000000000000",18104 => "0000000000000000",
18105 => "0000000000000000",18106 => "0000000000000000",
18107 => "0000000000000000",18108 => "0000000000000000",
18109 => "0000000000000000",18110 => "0000000000000000",
18111 => "0000000000000000",18112 => "0000000000000000",
18113 => "0000000000000000",18114 => "0000000000000000",
18115 => "0000000000000000",18116 => "0000000000000000",
18117 => "0000000000000000",18118 => "0000000000000000",
18119 => "0000000000000000",18120 => "0000000000000000",
18121 => "0000000000000000",18122 => "0000000000000000",
18123 => "0000000000000000",18124 => "0000000000000000",
18125 => "0000000000000000",18126 => "0000000000000000",
18127 => "0000000000000000",18128 => "0000000000000000",
18129 => "0000000000000000",18130 => "0000000000000000",
18131 => "0000000000000000",18132 => "0000000000000000",
18133 => "0000000000000000",18134 => "0000000000000000",
18135 => "0000000000000000",18136 => "0000000000000000",
18137 => "0000000000000000",18138 => "0000000000000000",
18139 => "0000000000000000",18140 => "0000000000000000",
18141 => "0000000000000000",18142 => "0000000000000000",
18143 => "0000000000000000",18144 => "0000000000000000",
18145 => "0000000000000000",18146 => "0000000000000000",
18147 => "0000000000000000",18148 => "0000000000000000",
18149 => "0000000000000000",18150 => "0000000000000000",
18151 => "0000000000000000",18152 => "0000000000000000",
18153 => "0000000000000000",18154 => "0000000000000000",
18155 => "0000000000000000",18156 => "0000000000000000",
18157 => "0000000000000000",18158 => "0000000000000000",
18159 => "0000000000000000",18160 => "0000000000000000",
18161 => "0000000000000000",18162 => "0000000000000000",
18163 => "0000000000000000",18164 => "0000000000000000",
18165 => "0000000000000000",18166 => "0000000000000000",
18167 => "0000000000000000",18168 => "0000000000000000",
18169 => "0000000000000000",18170 => "0000000000000000",
18171 => "0000000000000000",18172 => "0000000000000000",
18173 => "0000000000000000",18174 => "0000000000000000",
18175 => "0000000000000000",18176 => "0000000000000000",
18177 => "0000000000000000",18178 => "0000000000000000",
18179 => "0000000000000000",18180 => "0000000000000000",
18181 => "0000000000000000",18182 => "0000000000000000",
18183 => "0000000000000000",18184 => "0000000000000000",
18185 => "0000000000000000",18186 => "0000000000000000",
18187 => "0000000000000000",18188 => "0000000000000000",
18189 => "0000000000000000",18190 => "0000000000000000",
18191 => "0000000000000000",18192 => "0000000000000000",
18193 => "0000000000000000",18194 => "0000000000000000",
18195 => "0000000000000000",18196 => "0000000000000000",
18197 => "0000000000000000",18198 => "0000000000000000",
18199 => "0000000000000000",18200 => "0000000000000000",
18201 => "0000000000000000",18202 => "0000000000000000",
18203 => "0000000000000000",18204 => "0000000000000000",
18205 => "0000000000000000",18206 => "0000000000000000",
18207 => "0000000000000000",18208 => "0000000000000000",
18209 => "0000000000000000",18210 => "0000000000000000",
18211 => "0000000000000000",18212 => "0000000000000000",
18213 => "0000000000000000",18214 => "0000000000000000",
18215 => "0000000000000000",18216 => "0000000000000000",
18217 => "0000000000000000",18218 => "0000000000000000",
18219 => "0000000000000000",18220 => "0000000000000000",
18221 => "0000000000000000",18222 => "0000000000000000",
18223 => "0000000000000000",18224 => "0000000000000000",
18225 => "0000000000000000",18226 => "0000000000000000",
18227 => "0000000000000000",18228 => "0000000000000000",
18229 => "0000000000000000",18230 => "0000000000000000",
18231 => "0000000000000000",18232 => "0000000000000000",
18233 => "0000000000000000",18234 => "0000000000000000",
18235 => "0000000000000000",18236 => "0000000000000000",
18237 => "0000000000000000",18238 => "0000000000000000",
18239 => "0000000000000000",18240 => "0000000000000000",
18241 => "0000000000000000",18242 => "0000000000000000",
18243 => "0000000000000000",18244 => "0000000000000000",
18245 => "0000000000000000",18246 => "0000000000000000",
18247 => "0000000000000000",18248 => "0000000000000000",
18249 => "0000000000000000",18250 => "0000000000000000",
18251 => "0000000000000000",18252 => "0000000000000000",
18253 => "0000000000000000",18254 => "0000000000000000",
18255 => "0000000000000000",18256 => "0000000000000000",
18257 => "0000000000000000",18258 => "0000000000000000",
18259 => "0000000000000000",18260 => "0000000000000000",
18261 => "0000000000000000",18262 => "0000000000000000",
18263 => "0000000000000000",18264 => "0000000000000000",
18265 => "0000000000000000",18266 => "0000000000000000",
18267 => "0000000000000000",18268 => "0000000000000000",
18269 => "0000000000000000",18270 => "0000000000000000",
18271 => "0000000000000000",18272 => "0000000000000000",
18273 => "0000000000000000",18274 => "0000000000000000",
18275 => "0000000000000000",18276 => "0000000000000000",
18277 => "0000000000000000",18278 => "0000000000000000",
18279 => "0000000000000000",18280 => "0000000000000000",
18281 => "0000000000000000",18282 => "0000000000000000",
18283 => "0000000000000000",18284 => "0000000000000000",
18285 => "0000000000000000",18286 => "0000000000000000",
18287 => "0000000000000000",18288 => "0000000000000000",
18289 => "0000000000000000",18290 => "0000000000000000",
18291 => "0000000000000000",18292 => "0000000000000000",
18293 => "0000000000000000",18294 => "0000000000000000",
18295 => "0000000000000000",18296 => "0000000000000000",
18297 => "0000000000000000",18298 => "0000000000000000",
18299 => "0000000000000000",18300 => "0000000000000000",
18301 => "0000000000000000",18302 => "0000000000000000",
18303 => "0000000000000000",18304 => "0000000000000000",
18305 => "0000000000000000",18306 => "0000000000000000",
18307 => "0000000000000000",18308 => "0000000000000000",
18309 => "0000000000000000",18310 => "0000000000000000",
18311 => "0000000000000000",18312 => "0000000000000000",
18313 => "0000000000000000",18314 => "0000000000000000",
18315 => "0000000000000000",18316 => "0000000000000000",
18317 => "0000000000000000",18318 => "0000000000000000",
18319 => "0000000000000000",18320 => "0000000000000000",
18321 => "0000000000000000",18322 => "0000000000000000",
18323 => "0000000000000000",18324 => "0000000000000000",
18325 => "0000000000000000",18326 => "0000000000000000",
18327 => "0000000000000000",18328 => "0000000000000000",
18329 => "0000000000000000",18330 => "0000000000000000",
18331 => "0000000000000000",18332 => "0000000000000000",
18333 => "0000000000000000",18334 => "0000000000000000",
18335 => "0000000000000000",18336 => "0000000000000000",
18337 => "0000000000000000",18338 => "0000000000000000",
18339 => "0000000000000000",18340 => "0000000000000000",
18341 => "0000000000000000",18342 => "0000000000000000",
18343 => "0000000000000000",18344 => "0000000000000000",
18345 => "0000000000000000",18346 => "0000000000000000",
18347 => "0000000000000000",18348 => "0000000000000000",
18349 => "0000000000000000",18350 => "0000000000000000",
18351 => "0000000000000000",18352 => "0000000000000000",
18353 => "0000000000000000",18354 => "0000000000000000",
18355 => "0000000000000000",18356 => "0000000000000000",
18357 => "0000000000000000",18358 => "0000000000000000",
18359 => "0000000000000000",18360 => "0000000000000000",
18361 => "0000000000000000",18362 => "0000000000000000",
18363 => "0000000000000000",18364 => "0000000000000000",
18365 => "0000000000000000",18366 => "0000000000000000",
18367 => "0000000000000000",18368 => "0000000000000000",
18369 => "0000000000000000",18370 => "0000000000000000",
18371 => "0000000000000000",18372 => "0000000000000000",
18373 => "0000000000000000",18374 => "0000000000000000",
18375 => "0000000000000000",18376 => "0000000000000000",
18377 => "0000000000000000",18378 => "0000000000000000",
18379 => "0000000000000000",18380 => "0000000000000000",
18381 => "0000000000000000",18382 => "0000000000000000",
18383 => "0000000000000000",18384 => "0000000000000000",
18385 => "0000000000000000",18386 => "0000000000000000",
18387 => "0000000000000000",18388 => "0000000000000000",
18389 => "0000000000000000",18390 => "0000000000000000",
18391 => "0000000000000000",18392 => "0000000000000000",
18393 => "0000000000000000",18394 => "0000000000000000",
18395 => "0000000000000000",18396 => "0000000000000000",
18397 => "0000000000000000",18398 => "0000000000000000",
18399 => "0000000000000000",18400 => "0000000000000000",
18401 => "0000000000000000",18402 => "0000000000000000",
18403 => "0000000000000000",18404 => "0000000000000000",
18405 => "0000000000000000",18406 => "0000000000000000",
18407 => "0000000000000000",18408 => "0000000000000000",
18409 => "0000000000000000",18410 => "0000000000000000",
18411 => "0000000000000000",18412 => "0000000000000000",
18413 => "0000000000000000",18414 => "0000000000000000",
18415 => "0000000000000000",18416 => "0000000000000000",
18417 => "0000000000000000",18418 => "0000000000000000",
18419 => "0000000000000000",18420 => "0000000000000000",
18421 => "0000000000000000",18422 => "0000000000000000",
18423 => "0000000000000000",18424 => "0000000000000000",
18425 => "0000000000000000",18426 => "0000000000000000",
18427 => "0000000000000000",18428 => "0000000000000000",
18429 => "0000000000000000",18430 => "0000000000000000",
18431 => "0000000000000000",18432 => "0000000000000000",
18433 => "0000000000000000",18434 => "0000000000000000",
18435 => "0000000000000000",18436 => "0000000000000000",
18437 => "0000000000000000",18438 => "0000000000000000",
18439 => "0000000000000000",18440 => "0000000000000000",
18441 => "0000000000000000",18442 => "0000000000000000",
18443 => "0000000000000000",18444 => "0000000000000000",
18445 => "0000000000000000",18446 => "0000000000000000",
18447 => "0000000000000000",18448 => "0000000000000000",
18449 => "0000000000000000",18450 => "0000000000000000",
18451 => "0000000000000000",18452 => "0000000000000000",
18453 => "0000000000000000",18454 => "0000000000000000",
18455 => "0000000000000000",18456 => "0000000000000000",
18457 => "0000000000000000",18458 => "0000000000000000",
18459 => "0000000000000000",18460 => "0000000000000000",
18461 => "0000000000000000",18462 => "0000000000000000",
18463 => "0000000000000000",18464 => "0000000000000000",
18465 => "0000000000000000",18466 => "0000000000000000",
18467 => "0000000000000000",18468 => "0000000000000000",
18469 => "0000000000000000",18470 => "0000000000000000",
18471 => "0000000000000000",18472 => "0000000000000000",
18473 => "0000000000000000",18474 => "0000000000000000",
18475 => "0000000000000000",18476 => "0000000000000000",
18477 => "0000000000000000",18478 => "0000000000000000",
18479 => "0000000000000000",18480 => "0000000000000000",
18481 => "0000000000000000",18482 => "0000000000000000",
18483 => "0000000000000000",18484 => "0000000000000000",
18485 => "0000000000000000",18486 => "0000000000000000",
18487 => "0000000000000000",18488 => "0000000000000000",
18489 => "0000000000000000",18490 => "0000000000000000",
18491 => "0000000000000000",18492 => "0000000000000000",
18493 => "0000000000000000",18494 => "0000000000000000",
18495 => "0000000000000000",18496 => "0000000000000000",
18497 => "0000000000000000",18498 => "0000000000000000",
18499 => "0000000000000000",18500 => "0000000000000000",
18501 => "0000000000000000",18502 => "0000000000000000",
18503 => "0000000000000000",18504 => "0000000000000000",
18505 => "0000000000000000",18506 => "0000000000000000",
18507 => "0000000000000000",18508 => "0000000000000000",
18509 => "0000000000000000",18510 => "0000000000000000",
18511 => "0000000000000000",18512 => "0000000000000000",
18513 => "0000000000000000",18514 => "0000000000000000",
18515 => "0000000000000000",18516 => "0000000000000000",
18517 => "0000000000000000",18518 => "0000000000000000",
18519 => "0000000000000000",18520 => "0000000000000000",
18521 => "0000000000000000",18522 => "0000000000000000",
18523 => "0000000000000000",18524 => "0000000000000000",
18525 => "0000000000000000",18526 => "0000000000000000",
18527 => "0000000000000000",18528 => "0000000000000000",
18529 => "0000000000000000",18530 => "0000000000000000",
18531 => "0000000000000000",18532 => "0000000000000000",
18533 => "0000000000000000",18534 => "0000000000000000",
18535 => "0000000000000000",18536 => "0000000000000000",
18537 => "0000000000000000",18538 => "0000000000000000",
18539 => "0000000000000000",18540 => "0000000000000000",
18541 => "0000000000000000",18542 => "0000000000000000",
18543 => "0000000000000000",18544 => "0000000000000000",
18545 => "0000000000000000",18546 => "0000000000000000",
18547 => "0000000000000000",18548 => "0000000000000000",
18549 => "0000000000000000",18550 => "0000000000000000",
18551 => "0000000000000000",18552 => "0000000000000000",
18553 => "0000000000000000",18554 => "0000000000000000",
18555 => "0000000000000000",18556 => "0000000000000000",
18557 => "0000000000000000",18558 => "0000000000000000",
18559 => "0000000000000000",18560 => "0000000000000000",
18561 => "0000000000000000",18562 => "0000000000000000",
18563 => "0000000000000000",18564 => "0000000000000000",
18565 => "0000000000000000",18566 => "0000000000000000",
18567 => "0000000000000000",18568 => "0000000000000000",
18569 => "0000000000000000",18570 => "0000000000000000",
18571 => "0000000000000000",18572 => "0000000000000000",
18573 => "0000000000000000",18574 => "0000000000000000",
18575 => "0000000000000000",18576 => "0000000000000000",
18577 => "0000000000000000",18578 => "0000000000000000",
18579 => "0000000000000000",18580 => "0000000000000000",
18581 => "0000000000000000",18582 => "0000000000000000",
18583 => "0000000000000000",18584 => "0000000000000000",
18585 => "0000000000000000",18586 => "0000000000000000",
18587 => "0000000000000000",18588 => "0000000000000000",
18589 => "0000000000000000",18590 => "0000000000000000",
18591 => "0000000000000000",18592 => "0000000000000000",
18593 => "0000000000000000",18594 => "0000000000000000",
18595 => "0000000000000000",18596 => "0000000000000000",
18597 => "0000000000000000",18598 => "0000000000000000",
18599 => "0000000000000000",18600 => "0000000000000000",
18601 => "0000000000000000",18602 => "0000000000000000",
18603 => "0000000000000000",18604 => "0000000000000000",
18605 => "0000000000000000",18606 => "0000000000000000",
18607 => "0000000000000000",18608 => "0000000000000000",
18609 => "0000000000000000",18610 => "0000000000000000",
18611 => "0000000000000000",18612 => "0000000000000000",
18613 => "0000000000000000",18614 => "0000000000000000",
18615 => "0000000000000000",18616 => "0000000000000000",
18617 => "0000000000000000",18618 => "0000000000000000",
18619 => "0000000000000000",18620 => "0000000000000000",
18621 => "0000000000000000",18622 => "0000000000000000",
18623 => "0000000000000000",18624 => "0000000000000000",
18625 => "0000000000000000",18626 => "0000000000000000",
18627 => "0000000000000000",18628 => "0000000000000000",
18629 => "0000000000000000",18630 => "0000000000000000",
18631 => "0000000000000000",18632 => "0000000000000000",
18633 => "0000000000000000",18634 => "0000000000000000",
18635 => "0000000000000000",18636 => "0000000000000000",
18637 => "0000000000000000",18638 => "0000000000000000",
18639 => "0000000000000000",18640 => "0000000000000000",
18641 => "0000000000000000",18642 => "0000000000000000",
18643 => "0000000000000000",18644 => "0000000000000000",
18645 => "0000000000000000",18646 => "0000000000000000",
18647 => "0000000000000000",18648 => "0000000000000000",
18649 => "0000000000000000",18650 => "0000000000000000",
18651 => "0000000000000000",18652 => "0000000000000000",
18653 => "0000000000000000",18654 => "0000000000000000",
18655 => "0000000000000000",18656 => "0000000000000000",
18657 => "0000000000000000",18658 => "0000000000000000",
18659 => "0000000000000000",18660 => "0000000000000000",
18661 => "0000000000000000",18662 => "0000000000000000",
18663 => "0000000000000000",18664 => "0000000000000000",
18665 => "0000000000000000",18666 => "0000000000000000",
18667 => "0000000000000000",18668 => "0000000000000000",
18669 => "0000000000000000",18670 => "0000000000000000",
18671 => "0000000000000000",18672 => "0000000000000000",
18673 => "0000000000000000",18674 => "0000000000000000",
18675 => "0000000000000000",18676 => "0000000000000000",
18677 => "0000000000000000",18678 => "0000000000000000",
18679 => "0000000000000000",18680 => "0000000000000000",
18681 => "0000000000000000",18682 => "0000000000000000",
18683 => "0000000000000000",18684 => "0000000000000000",
18685 => "0000000000000000",18686 => "0000000000000000",
18687 => "0000000000000000",18688 => "0000000000000000",
18689 => "0000000000000000",18690 => "0000000000000000",
18691 => "0000000000000000",18692 => "0000000000000000",
18693 => "0000000000000000",18694 => "0000000000000000",
18695 => "0000000000000000",18696 => "0000000000000000",
18697 => "0000000000000000",18698 => "0000000000000000",
18699 => "0000000000000000",18700 => "0000000000000000",
18701 => "0000000000000000",18702 => "0000000000000000",
18703 => "0000000000000000",18704 => "0000000000000000",
18705 => "0000000000000000",18706 => "0000000000000000",
18707 => "0000000000000000",18708 => "0000000000000000",
18709 => "0000000000000000",18710 => "0000000000000000",
18711 => "0000000000000000",18712 => "0000000000000000",
18713 => "0000000000000000",18714 => "0000000000000000",
18715 => "0000000000000000",18716 => "0000000000000000",
18717 => "0000000000000000",18718 => "0000000000000000",
18719 => "0000000000000000",18720 => "0000000000000000",
18721 => "0000000000000000",18722 => "0000000000000000",
18723 => "0000000000000000",18724 => "0000000000000000",
18725 => "0000000000000000",18726 => "0000000000000000",
18727 => "0000000000000000",18728 => "0000000000000000",
18729 => "0000000000000000",18730 => "0000000000000000",
18731 => "0000000000000000",18732 => "0000000000000000",
18733 => "0000000000000000",18734 => "0000000000000000",
18735 => "0000000000000000",18736 => "0000000000000000",
18737 => "0000000000000000",18738 => "0000000000000000",
18739 => "0000000000000000",18740 => "0000000000000000",
18741 => "0000000000000000",18742 => "0000000000000000",
18743 => "0000000000000000",18744 => "0000000000000000",
18745 => "0000000000000000",18746 => "0000000000000000",
18747 => "0000000000000000",18748 => "0000000000000000",
18749 => "0000000000000000",18750 => "0000000000000000",
18751 => "0000000000000000",18752 => "0000000000000000",
18753 => "0000000000000000",18754 => "0000000000000000",
18755 => "0000000000000000",18756 => "0000000000000000",
18757 => "0000000000000000",18758 => "0000000000000000",
18759 => "0000000000000000",18760 => "0000000000000000",
18761 => "0000000000000000",18762 => "0000000000000000",
18763 => "0000000000000000",18764 => "0000000000000000",
18765 => "0000000000000000",18766 => "0000000000000000",
18767 => "0000000000000000",18768 => "0000000000000000",
18769 => "0000000000000000",18770 => "0000000000000000",
18771 => "0000000000000000",18772 => "0000000000000000",
18773 => "0000000000000000",18774 => "0000000000000000",
18775 => "0000000000000000",18776 => "0000000000000000",
18777 => "0000000000000000",18778 => "0000000000000000",
18779 => "0000000000000000",18780 => "0000000000000000",
18781 => "0000000000000000",18782 => "0000000000000000",
18783 => "0000000000000000",18784 => "0000000000000000",
18785 => "0000000000000000",18786 => "0000000000000000",
18787 => "0000000000000000",18788 => "0000000000000000",
18789 => "0000000000000000",18790 => "0000000000000000",
18791 => "0000000000000000",18792 => "0000000000000000",
18793 => "0000000000000000",18794 => "0000000000000000",
18795 => "0000000000000000",18796 => "0000000000000000",
18797 => "0000000000000000",18798 => "0000000000000000",
18799 => "0000000000000000",18800 => "0000000000000000",
18801 => "0000000000000000",18802 => "0000000000000000",
18803 => "0000000000000000",18804 => "0000000000000000",
18805 => "0000000000000000",18806 => "0000000000000000",
18807 => "0000000000000000",18808 => "0000000000000000",
18809 => "0000000000000000",18810 => "0000000000000000",
18811 => "0000000000000000",18812 => "0000000000000000",
18813 => "0000000000000000",18814 => "0000000000000000",
18815 => "0000000000000000",18816 => "0000000000000000",
18817 => "0000000000000000",18818 => "0000000000000000",
18819 => "0000000000000000",18820 => "0000000000000000",
18821 => "0000000000000000",18822 => "0000000000000000",
18823 => "0000000000000000",18824 => "0000000000000000",
18825 => "0000000000000000",18826 => "0000000000000000",
18827 => "0000000000000000",18828 => "0000000000000000",
18829 => "0000000000000000",18830 => "0000000000000000",
18831 => "0000000000000000",18832 => "0000000000000000",
18833 => "0000000000000000",18834 => "0000000000000000",
18835 => "0000000000000000",18836 => "0000000000000000",
18837 => "0000000000000000",18838 => "0000000000000000",
18839 => "0000000000000000",18840 => "0000000000000000",
18841 => "0000000000000000",18842 => "0000000000000000",
18843 => "0000000000000000",18844 => "0000000000000000",
18845 => "0000000000000000",18846 => "0000000000000000",
18847 => "0000000000000000",18848 => "0000000000000000",
18849 => "0000000000000000",18850 => "0000000000000000",
18851 => "0000000000000000",18852 => "0000000000000000",
18853 => "0000000000000000",18854 => "0000000000000000",
18855 => "0000000000000000",18856 => "0000000000000000",
18857 => "0000000000000000",18858 => "0000000000000000",
18859 => "0000000000000000",18860 => "0000000000000000",
18861 => "0000000000000000",18862 => "0000000000000000",
18863 => "0000000000000000",18864 => "0000000000000000",
18865 => "0000000000000000",18866 => "0000000000000000",
18867 => "0000000000000000",18868 => "0000000000000000",
18869 => "0000000000000000",18870 => "0000000000000000",
18871 => "0000000000000000",18872 => "0000000000000000",
18873 => "0000000000000000",18874 => "0000000000000000",
18875 => "0000000000000000",18876 => "0000000000000000",
18877 => "0000000000000000",18878 => "0000000000000000",
18879 => "0000000000000000",18880 => "0000000000000000",
18881 => "0000000000000000",18882 => "0000000000000000",
18883 => "0000000000000000",18884 => "0000000000000000",
18885 => "0000000000000000",18886 => "0000000000000000",
18887 => "0000000000000000",18888 => "0000000000000000",
18889 => "0000000000000000",18890 => "0000000000000000",
18891 => "0000000000000000",18892 => "0000000000000000",
18893 => "0000000000000000",18894 => "0000000000000000",
18895 => "0000000000000000",18896 => "0000000000000000",
18897 => "0000000000000000",18898 => "0000000000000000",
18899 => "0000000000000000",18900 => "0000000000000000",
18901 => "0000000000000000",18902 => "0000000000000000",
18903 => "0000000000000000",18904 => "0000000000000000",
18905 => "0000000000000000",18906 => "0000000000000000",
18907 => "0000000000000000",18908 => "0000000000000000",
18909 => "0000000000000000",18910 => "0000000000000000",
18911 => "0000000000000000",18912 => "0000000000000000",
18913 => "0000000000000000",18914 => "0000000000000000",
18915 => "0000000000000000",18916 => "0000000000000000",
18917 => "0000000000000000",18918 => "0000000000000000",
18919 => "0000000000000000",18920 => "0000000000000000",
18921 => "0000000000000000",18922 => "0000000000000000",
18923 => "0000000000000000",18924 => "0000000000000000",
18925 => "0000000000000000",18926 => "0000000000000000",
18927 => "0000000000000000",18928 => "0000000000000000",
18929 => "0000000000000000",18930 => "0000000000000000",
18931 => "0000000000000000",18932 => "0000000000000000",
18933 => "0000000000000000",18934 => "0000000000000000",
18935 => "0000000000000000",18936 => "0000000000000000",
18937 => "0000000000000000",18938 => "0000000000000000",
18939 => "0000000000000000",18940 => "0000000000000000",
18941 => "0000000000000000",18942 => "0000000000000000",
18943 => "0000000000000000",18944 => "0000000000000000",
18945 => "0000000000000000",18946 => "0000000000000000",
18947 => "0000000000000000",18948 => "0000000000000000",
18949 => "0000000000000000",18950 => "0000000000000000",
18951 => "0000000000000000",18952 => "0000000000000000",
18953 => "0000000000000000",18954 => "0000000000000000",
18955 => "0000000000000000",18956 => "0000000000000000",
18957 => "0000000000000000",18958 => "0000000000000000",
18959 => "0000000000000000",18960 => "0000000000000000",
18961 => "0000000000000000",18962 => "0000000000000000",
18963 => "0000000000000000",18964 => "0000000000000000",
18965 => "0000000000000000",18966 => "0000000000000000",
18967 => "0000000000000000",18968 => "0000000000000000",
18969 => "0000000000000000",18970 => "0000000000000000",
18971 => "0000000000000000",18972 => "0000000000000000",
18973 => "0000000000000000",18974 => "0000000000000000",
18975 => "0000000000000000",18976 => "0000000000000000",
18977 => "0000000000000000",18978 => "0000000000000000",
18979 => "0000000000000000",18980 => "0000000000000000",
18981 => "0000000000000000",18982 => "0000000000000000",
18983 => "0000000000000000",18984 => "0000000000000000",
18985 => "0000000000000000",18986 => "0000000000000000",
18987 => "0000000000000000",18988 => "0000000000000000",
18989 => "0000000000000000",18990 => "0000000000000000",
18991 => "0000000000000000",18992 => "0000000000000000",
18993 => "0000000000000000",18994 => "0000000000000000",
18995 => "0000000000000000",18996 => "0000000000000000",
18997 => "0000000000000000",18998 => "0000000000000000",
18999 => "0000000000000000",19000 => "0000000000000000",
19001 => "0000000000000000",19002 => "0000000000000000",
19003 => "0000000000000000",19004 => "0000000000000000",
19005 => "0000000000000000",19006 => "0000000000000000",
19007 => "0000000000000000",19008 => "0000000000000000",
19009 => "0000000000000000",19010 => "0000000000000000",
19011 => "0000000000000000",19012 => "0000000000000000",
19013 => "0000000000000000",19014 => "0000000000000000",
19015 => "0000000000000000",19016 => "0000000000000000",
19017 => "0000000000000000",19018 => "0000000000000000",
19019 => "0000000000000000",19020 => "0000000000000000",
19021 => "0000000000000000",19022 => "0000000000000000",
19023 => "0000000000000000",19024 => "0000000000000000",
19025 => "0000000000000000",19026 => "0000000000000000",
19027 => "0000000000000000",19028 => "0000000000000000",
19029 => "0000000000000000",19030 => "0000000000000000",
19031 => "0000000000000000",19032 => "0000000000000000",
19033 => "0000000000000000",19034 => "0000000000000000",
19035 => "0000000000000000",19036 => "0000000000000000",
19037 => "0000000000000000",19038 => "0000000000000000",
19039 => "0000000000000000",19040 => "0000000000000000",
19041 => "0000000000000000",19042 => "0000000000000000",
19043 => "0000000000000000",19044 => "0000000000000000",
19045 => "0000000000000000",19046 => "0000000000000000",
19047 => "0000000000000000",19048 => "0000000000000000",
19049 => "0000000000000000",19050 => "0000000000000000",
19051 => "0000000000000000",19052 => "0000000000000000",
19053 => "0000000000000000",19054 => "0000000000000000",
19055 => "0000000000000000",19056 => "0000000000000000",
19057 => "0000000000000000",19058 => "0000000000000000",
19059 => "0000000000000000",19060 => "0000000000000000",
19061 => "0000000000000000",19062 => "0000000000000000",
19063 => "0000000000000000",19064 => "0000000000000000",
19065 => "0000000000000000",19066 => "0000000000000000",
19067 => "0000000000000000",19068 => "0000000000000000",
19069 => "0000000000000000",19070 => "0000000000000000",
19071 => "0000000000000000",19072 => "0000000000000000",
19073 => "0000000000000000",19074 => "0000000000000000",
19075 => "0000000000000000",19076 => "0000000000000000",
19077 => "0000000000000000",19078 => "0000000000000000",
19079 => "0000000000000000",19080 => "0000000000000000",
19081 => "0000000000000000",19082 => "0000000000000000",
19083 => "0000000000000000",19084 => "0000000000000000",
19085 => "0000000000000000",19086 => "0000000000000000",
19087 => "0000000000000000",19088 => "0000000000000000",
19089 => "0000000000000000",19090 => "0000000000000000",
19091 => "0000000000000000",19092 => "0000000000000000",
19093 => "0000000000000000",19094 => "0000000000000000",
19095 => "0000000000000000",19096 => "0000000000000000",
19097 => "0000000000000000",19098 => "0000000000000000",
19099 => "0000000000000000",19100 => "0000000000000000",
19101 => "0000000000000000",19102 => "0000000000000000",
19103 => "0000000000000000",19104 => "0000000000000000",
19105 => "0000000000000000",19106 => "0000000000000000",
19107 => "0000000000000000",19108 => "0000000000000000",
19109 => "0000000000000000",19110 => "0000000000000000",
19111 => "0000000000000000",19112 => "0000000000000000",
19113 => "0000000000000000",19114 => "0000000000000000",
19115 => "0000000000000000",19116 => "0000000000000000",
19117 => "0000000000000000",19118 => "0000000000000000",
19119 => "0000000000000000",19120 => "0000000000000000",
19121 => "0000000000000000",19122 => "0000000000000000",
19123 => "0000000000000000",19124 => "0000000000000000",
19125 => "0000000000000000",19126 => "0000000000000000",
19127 => "0000000000000000",19128 => "0000000000000000",
19129 => "0000000000000000",19130 => "0000000000000000",
19131 => "0000000000000000",19132 => "0000000000000000",
19133 => "0000000000000000",19134 => "0000000000000000",
19135 => "0000000000000000",19136 => "0000000000000000",
19137 => "0000000000000000",19138 => "0000000000000000",
19139 => "0000000000000000",19140 => "0000000000000000",
19141 => "0000000000000000",19142 => "0000000000000000",
19143 => "0000000000000000",19144 => "0000000000000000",
19145 => "0000000000000000",19146 => "0000000000000000",
19147 => "0000000000000000",19148 => "0000000000000000",
19149 => "0000000000000000",19150 => "0000000000000000",
19151 => "0000000000000000",19152 => "0000000000000000",
19153 => "0000000000000000",19154 => "0000000000000000",
19155 => "0000000000000000",19156 => "0000000000000000",
19157 => "0000000000000000",19158 => "0000000000000000",
19159 => "0000000000000000",19160 => "0000000000000000",
19161 => "0000000000000000",19162 => "0000000000000000",
19163 => "0000000000000000",19164 => "0000000000000000",
19165 => "0000000000000000",19166 => "0000000000000000",
19167 => "0000000000000000",19168 => "0000000000000000",
19169 => "0000000000000000",19170 => "0000000000000000",
19171 => "0000000000000000",19172 => "0000000000000000",
19173 => "0000000000000000",19174 => "0000000000000000",
19175 => "0000000000000000",19176 => "0000000000000000",
19177 => "0000000000000000",19178 => "0000000000000000",
19179 => "0000000000000000",19180 => "0000000000000000",
19181 => "0000000000000000",19182 => "0000000000000000",
19183 => "0000000000000000",19184 => "0000000000000000",
19185 => "0000000000000000",19186 => "0000000000000000",
19187 => "0000000000000000",19188 => "0000000000000000",
19189 => "0000000000000000",19190 => "0000000000000000",
19191 => "0000000000000000",19192 => "0000000000000000",
19193 => "0000000000000000",19194 => "0000000000000000",
19195 => "0000000000000000",19196 => "0000000000000000",
19197 => "0000000000000000",19198 => "0000000000000000",
19199 => "0000000000000000",19200 => "0000000000000000",
19201 => "0000000000000000",19202 => "0000000000000000",
19203 => "0000000000000000",19204 => "0000000000000000",
19205 => "0000000000000000",19206 => "0000000000000000",
19207 => "0000000000000000",19208 => "0000000000000000",
19209 => "0000000000000000",19210 => "0000000000000000",
19211 => "0000000000000000",19212 => "0000000000000000",
19213 => "0000000000000000",19214 => "0000000000000000",
19215 => "0000000000000000",19216 => "0000000000000000",
19217 => "0000000000000000",19218 => "0000000000000000",
19219 => "0000000000000000",19220 => "0000000000000000",
19221 => "0000000000000000",19222 => "0000000000000000",
19223 => "0000000000000000",19224 => "0000000000000000",
19225 => "0000000000000000",19226 => "0000000000000000",
19227 => "0000000000000000",19228 => "0000000000000000",
19229 => "0000000000000000",19230 => "0000000000000000",
19231 => "0000000000000000",19232 => "0000000000000000",
19233 => "0000000000000000",19234 => "0000000000000000",
19235 => "0000000000000000",19236 => "0000000000000000",
19237 => "0000000000000000",19238 => "0000000000000000",
19239 => "0000000000000000",19240 => "0000000000000000",
19241 => "0000000000000000",19242 => "0000000000000000",
19243 => "0000000000000000",19244 => "0000000000000000",
19245 => "0000000000000000",19246 => "0000000000000000",
19247 => "0000000000000000",19248 => "0000000000000000",
19249 => "0000000000000000",19250 => "0000000000000000",
19251 => "0000000000000000",19252 => "0000000000000000",
19253 => "0000000000000000",19254 => "0000000000000000",
19255 => "0000000000000000",19256 => "0000000000000000",
19257 => "0000000000000000",19258 => "0000000000000000",
19259 => "0000000000000000",19260 => "0000000000000000",
19261 => "0000000000000000",19262 => "0000000000000000",
19263 => "0000000000000000",19264 => "0000000000000000",
19265 => "0000000000000000",19266 => "0000000000000000",
19267 => "0000000000000000",19268 => "0000000000000000",
19269 => "0000000000000000",19270 => "0000000000000000",
19271 => "0000000000000000",19272 => "0000000000000000",
19273 => "0000000000000000",19274 => "0000000000000000",
19275 => "0000000000000000",19276 => "0000000000000000",
19277 => "0000000000000000",19278 => "0000000000000000",
19279 => "0000000000000000",19280 => "0000000000000000",
19281 => "0000000000000000",19282 => "0000000000000000",
19283 => "0000000000000000",19284 => "0000000000000000",
19285 => "0000000000000000",19286 => "0000000000000000",
19287 => "0000000000000000",19288 => "0000000000000000",
19289 => "0000000000000000",19290 => "0000000000000000",
19291 => "0000000000000000",19292 => "0000000000000000",
19293 => "0000000000000000",19294 => "0000000000000000",
19295 => "0000000000000000",19296 => "0000000000000000",
19297 => "0000000000000000",19298 => "0000000000000000",
19299 => "0000000000000000",19300 => "0000000000000000",
19301 => "0000000000000000",19302 => "0000000000000000",
19303 => "0000000000000000",19304 => "0000000000000000",
19305 => "0000000000000000",19306 => "0000000000000000",
19307 => "0000000000000000",19308 => "0000000000000000",
19309 => "0000000000000000",19310 => "0000000000000000",
19311 => "0000000000000000",19312 => "0000000000000000",
19313 => "0000000000000000",19314 => "0000000000000000",
19315 => "0000000000000000",19316 => "0000000000000000",
19317 => "0000000000000000",19318 => "0000000000000000",
19319 => "0000000000000000",19320 => "0000000000000000",
19321 => "0000000000000000",19322 => "0000000000000000",
19323 => "0000000000000000",19324 => "0000000000000000",
19325 => "0000000000000000",19326 => "0000000000000000",
19327 => "0000000000000000",19328 => "0000000000000000",
19329 => "0000000000000000",19330 => "0000000000000000",
19331 => "0000000000000000",19332 => "0000000000000000",
19333 => "0000000000000000",19334 => "0000000000000000",
19335 => "0000000000000000",19336 => "0000000000000000",
19337 => "0000000000000000",19338 => "0000000000000000",
19339 => "0000000000000000",19340 => "0000000000000000",
19341 => "0000000000000000",19342 => "0000000000000000",
19343 => "0000000000000000",19344 => "0000000000000000",
19345 => "0000000000000000",19346 => "0000000000000000",
19347 => "0000000000000000",19348 => "0000000000000000",
19349 => "0000000000000000",19350 => "0000000000000000",
19351 => "0000000000000000",19352 => "0000000000000000",
19353 => "0000000000000000",19354 => "0000000000000000",
19355 => "0000000000000000",19356 => "0000000000000000",
19357 => "0000000000000000",19358 => "0000000000000000",
19359 => "0000000000000000",19360 => "0000000000000000",
19361 => "0000000000000000",19362 => "0000000000000000",
19363 => "0000000000000000",19364 => "0000000000000000",
19365 => "0000000000000000",19366 => "0000000000000000",
19367 => "0000000000000000",19368 => "0000000000000000",
19369 => "0000000000000000",19370 => "0000000000000000",
19371 => "0000000000000000",19372 => "0000000000000000",
19373 => "0000000000000000",19374 => "0000000000000000",
19375 => "0000000000000000",19376 => "0000000000000000",
19377 => "0000000000000000",19378 => "0000000000000000",
19379 => "0000000000000000",19380 => "0000000000000000",
19381 => "0000000000000000",19382 => "0000000000000000",
19383 => "0000000000000000",19384 => "0000000000000000",
19385 => "0000000000000000",19386 => "0000000000000000",
19387 => "0000000000000000",19388 => "0000000000000000",
19389 => "0000000000000000",19390 => "0000000000000000",
19391 => "0000000000000000",19392 => "0000000000000000",
19393 => "0000000000000000",19394 => "0000000000000000",
19395 => "0000000000000000",19396 => "0000000000000000",
19397 => "0000000000000000",19398 => "0000000000000000",
19399 => "0000000000000000",19400 => "0000000000000000",
19401 => "0000000000000000",19402 => "0000000000000000",
19403 => "0000000000000000",19404 => "0000000000000000",
19405 => "0000000000000000",19406 => "0000000000000000",
19407 => "0000000000000000",19408 => "0000000000000000",
19409 => "0000000000000000",19410 => "0000000000000000",
19411 => "0000000000000000",19412 => "0000000000000000",
19413 => "0000000000000000",19414 => "0000000000000000",
19415 => "0000000000000000",19416 => "0000000000000000",
19417 => "0000000000000000",19418 => "0000000000000000",
19419 => "0000000000000000",19420 => "0000000000000000",
19421 => "0000000000000000",19422 => "0000000000000000",
19423 => "0000000000000000",19424 => "0000000000000000",
19425 => "0000000000000000",19426 => "0000000000000000",
19427 => "0000000000000000",19428 => "0000000000000000",
19429 => "0000000000000000",19430 => "0000000000000000",
19431 => "0000000000000000",19432 => "0000000000000000",
19433 => "0000000000000000",19434 => "0000000000000000",
19435 => "0000000000000000",19436 => "0000000000000000",
19437 => "0000000000000000",19438 => "0000000000000000",
19439 => "0000000000000000",19440 => "0000000000000000",
19441 => "0000000000000000",19442 => "0000000000000000",
19443 => "0000000000000000",19444 => "0000000000000000",
19445 => "0000000000000000",19446 => "0000000000000000",
19447 => "0000000000000000",19448 => "0000000000000000",
19449 => "0000000000000000",19450 => "0000000000000000",
19451 => "0000000000000000",19452 => "0000000000000000",
19453 => "0000000000000000",19454 => "0000000000000000",
19455 => "0000000000000000",19456 => "0000000000000000",
19457 => "0000000000000000",19458 => "0000000000000000",
19459 => "0000000000000000",19460 => "0000000000000000",
19461 => "0000000000000000",19462 => "0000000000000000",
19463 => "0000000000000000",19464 => "0000000000000000",
19465 => "0000000000000000",19466 => "0000000000000000",
19467 => "0000000000000000",19468 => "0000000000000000",
19469 => "0000000000000000",19470 => "0000000000000000",
19471 => "0000000000000000",19472 => "0000000000000000",
19473 => "0000000000000000",19474 => "0000000000000000",
19475 => "0000000000000000",19476 => "0000000000000000",
19477 => "0000000000000000",19478 => "0000000000000000",
19479 => "0000000000000000",19480 => "0000000000000000",
19481 => "0000000000000000",19482 => "0000000000000000",
19483 => "0000000000000000",19484 => "0000000000000000",
19485 => "0000000000000000",19486 => "0000000000000000",
19487 => "0000000000000000",19488 => "0000000000000000",
19489 => "0000000000000000",19490 => "0000000000000000",
19491 => "0000000000000000",19492 => "0000000000000000",
19493 => "0000000000000000",19494 => "0000000000000000",
19495 => "0000000000000000",19496 => "0000000000000000",
19497 => "0000000000000000",19498 => "0000000000000000",
19499 => "0000000000000000",19500 => "0000000000000000",
19501 => "0000000000000000",19502 => "0000000000000000",
19503 => "0000000000000000",19504 => "0000000000000000",
19505 => "0000000000000000",19506 => "0000000000000000",
19507 => "0000000000000000",19508 => "0000000000000000",
19509 => "0000000000000000",19510 => "0000000000000000",
19511 => "0000000000000000",19512 => "0000000000000000",
19513 => "0000000000000000",19514 => "0000000000000000",
19515 => "0000000000000000",19516 => "0000000000000000",
19517 => "0000000000000000",19518 => "0000000000000000",
19519 => "0000000000000000",19520 => "0000000000000000",
19521 => "0000000000000000",19522 => "0000000000000000",
19523 => "0000000000000000",19524 => "0000000000000000",
19525 => "0000000000000000",19526 => "0000000000000000",
19527 => "0000000000000000",19528 => "0000000000000000",
19529 => "0000000000000000",19530 => "0000000000000000",
19531 => "0000000000000000",19532 => "0000000000000000",
19533 => "0000000000000000",19534 => "0000000000000000",
19535 => "0000000000000000",19536 => "0000000000000000",
19537 => "0000000000000000",19538 => "0000000000000000",
19539 => "0000000000000000",19540 => "0000000000000000",
19541 => "0000000000000000",19542 => "0000000000000000",
19543 => "0000000000000000",19544 => "0000000000000000",
19545 => "0000000000000000",19546 => "0000000000000000",
19547 => "0000000000000000",19548 => "0000000000000000",
19549 => "0000000000000000",19550 => "0000000000000000",
19551 => "0000000000000000",19552 => "0000000000000000",
19553 => "0000000000000000",19554 => "0000000000000000",
19555 => "0000000000000000",19556 => "0000000000000000",
19557 => "0000000000000000",19558 => "0000000000000000",
19559 => "0000000000000000",19560 => "0000000000000000",
19561 => "0000000000000000",19562 => "0000000000000000",
19563 => "0000000000000000",19564 => "0000000000000000",
19565 => "0000000000000000",19566 => "0000000000000000",
19567 => "0000000000000000",19568 => "0000000000000000",
19569 => "0000000000000000",19570 => "0000000000000000",
19571 => "0000000000000000",19572 => "0000000000000000",
19573 => "0000000000000000",19574 => "0000000000000000",
19575 => "0000000000000000",19576 => "0000000000000000",
19577 => "0000000000000000",19578 => "0000000000000000",
19579 => "0000000000000000",19580 => "0000000000000000",
19581 => "0000000000000000",19582 => "0000000000000000",
19583 => "0000000000000000",19584 => "0000000000000000",
19585 => "0000000000000000",19586 => "0000000000000000",
19587 => "0000000000000000",19588 => "0000000000000000",
19589 => "0000000000000000",19590 => "0000000000000000",
19591 => "0000000000000000",19592 => "0000000000000000",
19593 => "0000000000000000",19594 => "0000000000000000",
19595 => "0000000000000000",19596 => "0000000000000000",
19597 => "0000000000000000",19598 => "0000000000000000",
19599 => "0000000000000000",19600 => "0000000000000000",
19601 => "0000000000000000",19602 => "0000000000000000",
19603 => "0000000000000000",19604 => "0000000000000000",
19605 => "0000000000000000",19606 => "0000000000000000",
19607 => "0000000000000000",19608 => "0000000000000000",
19609 => "0000000000000000",19610 => "0000000000000000",
19611 => "0000000000000000",19612 => "0000000000000000",
19613 => "0000000000000000",19614 => "0000000000000000",
19615 => "0000000000000000",19616 => "0000000000000000",
19617 => "0000000000000000",19618 => "0000000000000000",
19619 => "0000000000000000",19620 => "0000000000000000",
19621 => "0000000000000000",19622 => "0000000000000000",
19623 => "0000000000000000",19624 => "0000000000000000",
19625 => "0000000000000000",19626 => "0000000000000000",
19627 => "0000000000000000",19628 => "0000000000000000",
19629 => "0000000000000000",19630 => "0000000000000000",
19631 => "0000000000000000",19632 => "0000000000000000",
19633 => "0000000000000000",19634 => "0000000000000000",
19635 => "0000000000000000",19636 => "0000000000000000",
19637 => "0000000000000000",19638 => "0000000000000000",
19639 => "0000000000000000",19640 => "0000000000000000",
19641 => "0000000000000000",19642 => "0000000000000000",
19643 => "0000000000000000",19644 => "0000000000000000",
19645 => "0000000000000000",19646 => "0000000000000000",
19647 => "0000000000000000",19648 => "0000000000000000",
19649 => "0000000000000000",19650 => "0000000000000000",
19651 => "0000000000000000",19652 => "0000000000000000",
19653 => "0000000000000000",19654 => "0000000000000000",
19655 => "0000000000000000",19656 => "0000000000000000",
19657 => "0000000000000000",19658 => "0000000000000000",
19659 => "0000000000000000",19660 => "0000000000000000",
19661 => "0000000000000000",19662 => "0000000000000000",
19663 => "0000000000000000",19664 => "0000000000000000",
19665 => "0000000000000000",19666 => "0000000000000000",
19667 => "0000000000000000",19668 => "0000000000000000",
19669 => "0000000000000000",19670 => "0000000000000000",
19671 => "0000000000000000",19672 => "0000000000000000",
19673 => "0000000000000000",19674 => "0000000000000000",
19675 => "0000000000000000",19676 => "0000000000000000",
19677 => "0000000000000000",19678 => "0000000000000000",
19679 => "0000000000000000",19680 => "0000000000000000",
19681 => "0000000000000000",19682 => "0000000000000000",
19683 => "0000000000000000",19684 => "0000000000000000",
19685 => "0000000000000000",19686 => "0000000000000000",
19687 => "0000000000000000",19688 => "0000000000000000",
19689 => "0000000000000000",19690 => "0000000000000000",
19691 => "0000000000000000",19692 => "0000000000000000",
19693 => "0000000000000000",19694 => "0000000000000000",
19695 => "0000000000000000",19696 => "0000000000000000",
19697 => "0000000000000000",19698 => "0000000000000000",
19699 => "0000000000000000",19700 => "0000000000000000",
19701 => "0000000000000000",19702 => "0000000000000000",
19703 => "0000000000000000",19704 => "0000000000000000",
19705 => "0000000000000000",19706 => "0000000000000000",
19707 => "0000000000000000",19708 => "0000000000000000",
19709 => "0000000000000000",19710 => "0000000000000000",
19711 => "0000000000000000",19712 => "0000000000000000",
19713 => "0000000000000000",19714 => "0000000000000000",
19715 => "0000000000000000",19716 => "0000000000000000",
19717 => "0000000000000000",19718 => "0000000000000000",
19719 => "0000000000000000",19720 => "0000000000000000",
19721 => "0000000000000000",19722 => "0000000000000000",
19723 => "0000000000000000",19724 => "0000000000000000",
19725 => "0000000000000000",19726 => "0000000000000000",
19727 => "0000000000000000",19728 => "0000000000000000",
19729 => "0000000000000000",19730 => "0000000000000000",
19731 => "0000000000000000",19732 => "0000000000000000",
19733 => "0000000000000000",19734 => "0000000000000000",
19735 => "0000000000000000",19736 => "0000000000000000",
19737 => "0000000000000000",19738 => "0000000000000000",
19739 => "0000000000000000",19740 => "0000000000000000",
19741 => "0000000000000000",19742 => "0000000000000000",
19743 => "0000000000000000",19744 => "0000000000000000",
19745 => "0000000000000000",19746 => "0000000000000000",
19747 => "0000000000000000",19748 => "0000000000000000",
19749 => "0000000000000000",19750 => "0000000000000000",
19751 => "0000000000000000",19752 => "0000000000000000",
19753 => "0000000000000000",19754 => "0000000000000000",
19755 => "0000000000000000",19756 => "0000000000000000",
19757 => "0000000000000000",19758 => "0000000000000000",
19759 => "0000000000000000",19760 => "0000000000000000",
19761 => "0000000000000000",19762 => "0000000000000000",
19763 => "0000000000000000",19764 => "0000000000000000",
19765 => "0000000000000000",19766 => "0000000000000000",
19767 => "0000000000000000",19768 => "0000000000000000",
19769 => "0000000000000000",19770 => "0000000000000000",
19771 => "0000000000000000",19772 => "0000000000000000",
19773 => "0000000000000000",19774 => "0000000000000000",
19775 => "0000000000000000",19776 => "0000000000000000",
19777 => "0000000000000000",19778 => "0000000000000000",
19779 => "0000000000000000",19780 => "0000000000000000",
19781 => "0000000000000000",19782 => "0000000000000000",
19783 => "0000000000000000",19784 => "0000000000000000",
19785 => "0000000000000000",19786 => "0000000000000000",
19787 => "0000000000000000",19788 => "0000000000000000",
19789 => "0000000000000000",19790 => "0000000000000000",
19791 => "0000000000000000",19792 => "0000000000000000",
19793 => "0000000000000000",19794 => "0000000000000000",
19795 => "0000000000000000",19796 => "0000000000000000",
19797 => "0000000000000000",19798 => "0000000000000000",
19799 => "0000000000000000",19800 => "0000000000000000",
19801 => "0000000000000000",19802 => "0000000000000000",
19803 => "0000000000000000",19804 => "0000000000000000",
19805 => "0000000000000000",19806 => "0000000000000000",
19807 => "0000000000000000",19808 => "0000000000000000",
19809 => "0000000000000000",19810 => "0000000000000000",
19811 => "0000000000000000",19812 => "0000000000000000",
19813 => "0000000000000000",19814 => "0000000000000000",
19815 => "0000000000000000",19816 => "0000000000000000",
19817 => "0000000000000000",19818 => "0000000000000000",
19819 => "0000000000000000",19820 => "0000000000000000",
19821 => "0000000000000000",19822 => "0000000000000000",
19823 => "0000000000000000",19824 => "0000000000000000",
19825 => "0000000000000000",19826 => "0000000000000000",
19827 => "0000000000000000",19828 => "0000000000000000",
19829 => "0000000000000000",19830 => "0000000000000000",
19831 => "0000000000000000",19832 => "0000000000000000",
19833 => "0000000000000000",19834 => "0000000000000000",
19835 => "0000000000000000",19836 => "0000000000000000",
19837 => "0000000000000000",19838 => "0000000000000000",
19839 => "0000000000000000",19840 => "0000000000000000",
19841 => "0000000000000000",19842 => "0000000000000000",
19843 => "0000000000000000",19844 => "0000000000000000",
19845 => "0000000000000000",19846 => "0000000000000000",
19847 => "0000000000000000",19848 => "0000000000000000",
19849 => "0000000000000000",19850 => "0000000000000000",
19851 => "0000000000000000",19852 => "0000000000000000",
19853 => "0000000000000000",19854 => "0000000000000000",
19855 => "0000000000000000",19856 => "0000000000000000",
19857 => "0000000000000000",19858 => "0000000000000000",
19859 => "0000000000000000",19860 => "0000000000000000",
19861 => "0000000000000000",19862 => "0000000000000000",
19863 => "0000000000000000",19864 => "0000000000000000",
19865 => "0000000000000000",19866 => "0000000000000000",
19867 => "0000000000000000",19868 => "0000000000000000",
19869 => "0000000000000000",19870 => "0000000000000000",
19871 => "0000000000000000",19872 => "0000000000000000",
19873 => "0000000000000000",19874 => "0000000000000000",
19875 => "0000000000000000",19876 => "0000000000000000",
19877 => "0000000000000000",19878 => "0000000000000000",
19879 => "0000000000000000",19880 => "0000000000000000",
19881 => "0000000000000000",19882 => "0000000000000000",
19883 => "0000000000000000",19884 => "0000000000000000",
19885 => "0000000000000000",19886 => "0000000000000000",
19887 => "0000000000000000",19888 => "0000000000000000",
19889 => "0000000000000000",19890 => "0000000000000000",
19891 => "0000000000000000",19892 => "0000000000000000",
19893 => "0000000000000000",19894 => "0000000000000000",
19895 => "0000000000000000",19896 => "0000000000000000",
19897 => "0000000000000000",19898 => "0000000000000000",
19899 => "0000000000000000",19900 => "0000000000000000",
19901 => "0000000000000000",19902 => "0000000000000000",
19903 => "0000000000000000",19904 => "0000000000000000",
19905 => "0000000000000000",19906 => "0000000000000000",
19907 => "0000000000000000",19908 => "0000000000000000",
19909 => "0000000000000000",19910 => "0000000000000000",
19911 => "0000000000000000",19912 => "0000000000000000",
19913 => "0000000000000000",19914 => "0000000000000000",
19915 => "0000000000000000",19916 => "0000000000000000",
19917 => "0000000000000000",19918 => "0000000000000000",
19919 => "0000000000000000",19920 => "0000000000000000",
19921 => "0000000000000000",19922 => "0000000000000000",
19923 => "0000000000000000",19924 => "0000000000000000",
19925 => "0000000000000000",19926 => "0000000000000000",
19927 => "0000000000000000",19928 => "0000000000000000",
19929 => "0000000000000000",19930 => "0000000000000000",
19931 => "0000000000000000",19932 => "0000000000000000",
19933 => "0000000000000000",19934 => "0000000000000000",
19935 => "0000000000000000",19936 => "0000000000000000",
19937 => "0000000000000000",19938 => "0000000000000000",
19939 => "0000000000000000",19940 => "0000000000000000",
19941 => "0000000000000000",19942 => "0000000000000000",
19943 => "0000000000000000",19944 => "0000000000000000",
19945 => "0000000000000000",19946 => "0000000000000000",
19947 => "0000000000000000",19948 => "0000000000000000",
19949 => "0000000000000000",19950 => "0000000000000000",
19951 => "0000000000000000",19952 => "0000000000000000",
19953 => "0000000000000000",19954 => "0000000000000000",
19955 => "0000000000000000",19956 => "0000000000000000",
19957 => "0000000000000000",19958 => "0000000000000000",
19959 => "0000000000000000",19960 => "0000000000000000",
19961 => "0000000000000000",19962 => "0000000000000000",
19963 => "0000000000000000",19964 => "0000000000000000",
19965 => "0000000000000000",19966 => "0000000000000000",
19967 => "0000000000000000",19968 => "0000000000000000",
19969 => "0000000000000000",19970 => "0000000000000000",
19971 => "0000000000000000",19972 => "0000000000000000",
19973 => "0000000000000000",19974 => "0000000000000000",
19975 => "0000000000000000",19976 => "0000000000000000",
19977 => "0000000000000000",19978 => "0000000000000000",
19979 => "0000000000000000",19980 => "0000000000000000",
19981 => "0000000000000000",19982 => "0000000000000000",
19983 => "0000000000000000",19984 => "0000000000000000",
19985 => "0000000000000000",19986 => "0000000000000000",
19987 => "0000000000000000",19988 => "0000000000000000",
19989 => "0000000000000000",19990 => "0000000000000000",
19991 => "0000000000000000",19992 => "0000000000000000",
19993 => "0000000000000000",19994 => "0000000000000000",
19995 => "0000000000000000",19996 => "0000000000000000",
19997 => "0000000000000000",19998 => "0000000000000000",
19999 => "0000000000000000",20000 => "0000000000000000",
20001 => "0000000000000000",20002 => "0000000000000000",
20003 => "0000000000000000",20004 => "0000000000000000",
20005 => "0000000000000000",20006 => "0000000000000000",
20007 => "0000000000000000",20008 => "0000000000000000",
20009 => "0000000000000000",20010 => "0000000000000000",
20011 => "0000000000000000",20012 => "0000000000000000",
20013 => "0000000000000000",20014 => "0000000000000000",
20015 => "0000000000000000",20016 => "0000000000000000",
20017 => "0000000000000000",20018 => "0000000000000000",
20019 => "0000000000000000",20020 => "0000000000000000",
20021 => "0000000000000000",20022 => "0000000000000000",
20023 => "0000000000000000",20024 => "0000000000000000",
20025 => "0000000000000000",20026 => "0000000000000000",
20027 => "0000000000000000",20028 => "0000000000000000",
20029 => "0000000000000000",20030 => "0000000000000000",
20031 => "0000000000000000",20032 => "0000000000000000",
20033 => "0000000000000000",20034 => "0000000000000000",
20035 => "0000000000000000",20036 => "0000000000000000",
20037 => "0000000000000000",20038 => "0000000000000000",
20039 => "0000000000000000",20040 => "0000000000000000",
20041 => "0000000000000000",20042 => "0000000000000000",
20043 => "0000000000000000",20044 => "0000000000000000",
20045 => "0000000000000000",20046 => "0000000000000000",
20047 => "0000000000000000",20048 => "0000000000000000",
20049 => "0000000000000000",20050 => "0000000000000000",
20051 => "0000000000000000",20052 => "0000000000000000",
20053 => "0000000000000000",20054 => "0000000000000000",
20055 => "0000000000000000",20056 => "0000000000000000",
20057 => "0000000000000000",20058 => "0000000000000000",
20059 => "0000000000000000",20060 => "0000000000000000",
20061 => "0000000000000000",20062 => "0000000000000000",
20063 => "0000000000000000",20064 => "0000000000000000",
20065 => "0000000000000000",20066 => "0000000000000000",
20067 => "0000000000000000",20068 => "0000000000000000",
20069 => "0000000000000000",20070 => "0000000000000000",
20071 => "0000000000000000",20072 => "0000000000000000",
20073 => "0000000000000000",20074 => "0000000000000000",
20075 => "0000000000000000",20076 => "0000000000000000",
20077 => "0000000000000000",20078 => "0000000000000000",
20079 => "0000000000000000",20080 => "0000000000000000",
20081 => "0000000000000000",20082 => "0000000000000000",
20083 => "0000000000000000",20084 => "0000000000000000",
20085 => "0000000000000000",20086 => "0000000000000000",
20087 => "0000000000000000",20088 => "0000000000000000",
20089 => "0000000000000000",20090 => "0000000000000000",
20091 => "0000000000000000",20092 => "0000000000000000",
20093 => "0000000000000000",20094 => "0000000000000000",
20095 => "0000000000000000",20096 => "0000000000000000",
20097 => "0000000000000000",20098 => "0000000000000000",
20099 => "0000000000000000",20100 => "0000000000000000",
20101 => "0000000000000000",20102 => "0000000000000000",
20103 => "0000000000000000",20104 => "0000000000000000",
20105 => "0000000000000000",20106 => "0000000000000000",
20107 => "0000000000000000",20108 => "0000000000000000",
20109 => "0000000000000000",20110 => "0000000000000000",
20111 => "0000000000000000",20112 => "0000000000000000",
20113 => "0000000000000000",20114 => "0000000000000000",
20115 => "0000000000000000",20116 => "0000000000000000",
20117 => "0000000000000000",20118 => "0000000000000000",
20119 => "0000000000000000",20120 => "0000000000000000",
20121 => "0000000000000000",20122 => "0000000000000000",
20123 => "0000000000000000",20124 => "0000000000000000",
20125 => "0000000000000000",20126 => "0000000000000000",
20127 => "0000000000000000",20128 => "0000000000000000",
20129 => "0000000000000000",20130 => "0000000000000000",
20131 => "0000000000000000",20132 => "0000000000000000",
20133 => "0000000000000000",20134 => "0000000000000000",
20135 => "0000000000000000",20136 => "0000000000000000",
20137 => "0000000000000000",20138 => "0000000000000000",
20139 => "0000000000000000",20140 => "0000000000000000",
20141 => "0000000000000000",20142 => "0000000000000000",
20143 => "0000000000000000",20144 => "0000000000000000",
20145 => "0000000000000000",20146 => "0000000000000000",
20147 => "0000000000000000",20148 => "0000000000000000",
20149 => "0000000000000000",20150 => "0000000000000000",
20151 => "0000000000000000",20152 => "0000000000000000",
20153 => "0000000000000000",20154 => "0000000000000000",
20155 => "0000000000000000",20156 => "0000000000000000",
20157 => "0000000000000000",20158 => "0000000000000000",
20159 => "0000000000000000",20160 => "0000000000000000",
20161 => "0000000000000000",20162 => "0000000000000000",
20163 => "0000000000000000",20164 => "0000000000000000",
20165 => "0000000000000000",20166 => "0000000000000000",
20167 => "0000000000000000",20168 => "0000000000000000",
20169 => "0000000000000000",20170 => "0000000000000000",
20171 => "0000000000000000",20172 => "0000000000000000",
20173 => "0000000000000000",20174 => "0000000000000000",
20175 => "0000000000000000",20176 => "0000000000000000",
20177 => "0000000000000000",20178 => "0000000000000000",
20179 => "0000000000000000",20180 => "0000000000000000",
20181 => "0000000000000000",20182 => "0000000000000000",
20183 => "0000000000000000",20184 => "0000000000000000",
20185 => "0000000000000000",20186 => "0000000000000000",
20187 => "0000000000000000",20188 => "0000000000000000",
20189 => "0000000000000000",20190 => "0000000000000000",
20191 => "0000000000000000",20192 => "0000000000000000",
20193 => "0000000000000000",20194 => "0000000000000000",
20195 => "0000000000000000",20196 => "0000000000000000",
20197 => "0000000000000000",20198 => "0000000000000000",
20199 => "0000000000000000",20200 => "0000000000000000",
20201 => "0000000000000000",20202 => "0000000000000000",
20203 => "0000000000000000",20204 => "0000000000000000",
20205 => "0000000000000000",20206 => "0000000000000000",
20207 => "0000000000000000",20208 => "0000000000000000",
20209 => "0000000000000000",20210 => "0000000000000000",
20211 => "0000000000000000",20212 => "0000000000000000",
20213 => "0000000000000000",20214 => "0000000000000000",
20215 => "0000000000000000",20216 => "0000000000000000",
20217 => "0000000000000000",20218 => "0000000000000000",
20219 => "0000000000000000",20220 => "0000000000000000",
20221 => "0000000000000000",20222 => "0000000000000000",
20223 => "0000000000000000",20224 => "0000000000000000",
20225 => "0000000000000000",20226 => "0000000000000000",
20227 => "0000000000000000",20228 => "0000000000000000",
20229 => "0000000000000000",20230 => "0000000000000000",
20231 => "0000000000000000",20232 => "0000000000000000",
20233 => "0000000000000000",20234 => "0000000000000000",
20235 => "0000000000000000",20236 => "0000000000000000",
20237 => "0000000000000000",20238 => "0000000000000000",
20239 => "0000000000000000",20240 => "0000000000000000",
20241 => "0000000000000000",20242 => "0000000000000000",
20243 => "0000000000000000",20244 => "0000000000000000",
20245 => "0000000000000000",20246 => "0000000000000000",
20247 => "0000000000000000",20248 => "0000000000000000",
20249 => "0000000000000000",20250 => "0000000000000000",
20251 => "0000000000000000",20252 => "0000000000000000",
20253 => "0000000000000000",20254 => "0000000000000000",
20255 => "0000000000000000",20256 => "0000000000000000",
20257 => "0000000000000000",20258 => "0000000000000000",
20259 => "0000000000000000",20260 => "0000000000000000",
20261 => "0000000000000000",20262 => "0000000000000000",
20263 => "0000000000000000",20264 => "0000000000000000",
20265 => "0000000000000000",20266 => "0000000000000000",
20267 => "0000000000000000",20268 => "0000000000000000",
20269 => "0000000000000000",20270 => "0000000000000000",
20271 => "0000000000000000",20272 => "0000000000000000",
20273 => "0000000000000000",20274 => "0000000000000000",
20275 => "0000000000000000",20276 => "0000000000000000",
20277 => "0000000000000000",20278 => "0000000000000000",
20279 => "0000000000000000",20280 => "0000000000000000",
20281 => "0000000000000000",20282 => "0000000000000000",
20283 => "0000000000000000",20284 => "0000000000000000",
20285 => "0000000000000000",20286 => "0000000000000000",
20287 => "0000000000000000",20288 => "0000000000000000",
20289 => "0000000000000000",20290 => "0000000000000000",
20291 => "0000000000000000",20292 => "0000000000000000",
20293 => "0000000000000000",20294 => "0000000000000000",
20295 => "0000000000000000",20296 => "0000000000000000",
20297 => "0000000000000000",20298 => "0000000000000000",
20299 => "0000000000000000",20300 => "0000000000000000",
20301 => "0000000000000000",20302 => "0000000000000000",
20303 => "0000000000000000",20304 => "0000000000000000",
20305 => "0000000000000000",20306 => "0000000000000000",
20307 => "0000000000000000",20308 => "0000000000000000",
20309 => "0000000000000000",20310 => "0000000000000000",
20311 => "0000000000000000",20312 => "0000000000000000",
20313 => "0000000000000000",20314 => "0000000000000000",
20315 => "0000000000000000",20316 => "0000000000000000",
20317 => "0000000000000000",20318 => "0000000000000000",
20319 => "0000000000000000",20320 => "0000000000000000",
20321 => "0000000000000000",20322 => "0000000000000000",
20323 => "0000000000000000",20324 => "0000000000000000",
20325 => "0000000000000000",20326 => "0000000000000000",
20327 => "0000000000000000",20328 => "0000000000000000",
20329 => "0000000000000000",20330 => "0000000000000000",
20331 => "0000000000000000",20332 => "0000000000000000",
20333 => "0000000000000000",20334 => "0000000000000000",
20335 => "0000000000000000",20336 => "0000000000000000",
20337 => "0000000000000000",20338 => "0000000000000000",
20339 => "0000000000000000",20340 => "0000000000000000",
20341 => "0000000000000000",20342 => "0000000000000000",
20343 => "0000000000000000",20344 => "0000000000000000",
20345 => "0000000000000000",20346 => "0000000000000000",
20347 => "0000000000000000",20348 => "0000000000000000",
20349 => "0000000000000000",20350 => "0000000000000000",
20351 => "0000000000000000",20352 => "0000000000000000",
20353 => "0000000000000000",20354 => "0000000000000000",
20355 => "0000000000000000",20356 => "0000000000000000",
20357 => "0000000000000000",20358 => "0000000000000000",
20359 => "0000000000000000",20360 => "0000000000000000",
20361 => "0000000000000000",20362 => "0000000000000000",
20363 => "0000000000000000",20364 => "0000000000000000",
20365 => "0000000000000000",20366 => "0000000000000000",
20367 => "0000000000000000",20368 => "0000000000000000",
20369 => "0000000000000000",20370 => "0000000000000000",
20371 => "0000000000000000",20372 => "0000000000000000",
20373 => "0000000000000000",20374 => "0000000000000000",
20375 => "0000000000000000",20376 => "0000000000000000",
20377 => "0000000000000000",20378 => "0000000000000000",
20379 => "0000000000000000",20380 => "0000000000000000",
20381 => "0000000000000000",20382 => "0000000000000000",
20383 => "0000000000000000",20384 => "0000000000000000",
20385 => "0000000000000000",20386 => "0000000000000000",
20387 => "0000000000000000",20388 => "0000000000000000",
20389 => "0000000000000000",20390 => "0000000000000000",
20391 => "0000000000000000",20392 => "0000000000000000",
20393 => "0000000000000000",20394 => "0000000000000000",
20395 => "0000000000000000",20396 => "0000000000000000",
20397 => "0000000000000000",20398 => "0000000000000000",
20399 => "0000000000000000",20400 => "0000000000000000",
20401 => "0000000000000000",20402 => "0000000000000000",
20403 => "0000000000000000",20404 => "0000000000000000",
20405 => "0000000000000000",20406 => "0000000000000000",
20407 => "0000000000000000",20408 => "0000000000000000",
20409 => "0000000000000000",20410 => "0000000000000000",
20411 => "0000000000000000",20412 => "0000000000000000",
20413 => "0000000000000000",20414 => "0000000000000000",
20415 => "0000000000000000",20416 => "0000000000000000",
20417 => "0000000000000000",20418 => "0000000000000000",
20419 => "0000000000000000",20420 => "0000000000000000",
20421 => "0000000000000000",20422 => "0000000000000000",
20423 => "0000000000000000",20424 => "0000000000000000",
20425 => "0000000000000000",20426 => "0000000000000000",
20427 => "0000000000000000",20428 => "0000000000000000",
20429 => "0000000000000000",20430 => "0000000000000000",
20431 => "0000000000000000",20432 => "0000000000000000",
20433 => "0000000000000000",20434 => "0000000000000000",
20435 => "0000000000000000",20436 => "0000000000000000",
20437 => "0000000000000000",20438 => "0000000000000000",
20439 => "0000000000000000",20440 => "0000000000000000",
20441 => "0000000000000000",20442 => "0000000000000000",
20443 => "0000000000000000",20444 => "0000000000000000",
20445 => "0000000000000000",20446 => "0000000000000000",
20447 => "0000000000000000",20448 => "0000000000000000",
20449 => "0000000000000000",20450 => "0000000000000000",
20451 => "0000000000000000",20452 => "0000000000000000",
20453 => "0000000000000000",20454 => "0000000000000000",
20455 => "0000000000000000",20456 => "0000000000000000",
20457 => "0000000000000000",20458 => "0000000000000000",
20459 => "0000000000000000",20460 => "0000000000000000",
20461 => "0000000000000000",20462 => "0000000000000000",
20463 => "0000000000000000",20464 => "0000000000000000",
20465 => "0000000000000000",20466 => "0000000000000000",
20467 => "0000000000000000",20468 => "0000000000000000",
20469 => "0000000000000000",20470 => "0000000000000000",
20471 => "0000000000000000",20472 => "0000000000000000",
20473 => "0000000000000000",20474 => "0000000000000000",
20475 => "0000000000000000",20476 => "0000000000000000",
20477 => "0000000000000000",20478 => "0000000000000000",
20479 => "0000000000000000",20480 => "0000000000000000",
20481 => "0000000000000000",20482 => "0000000000000000",
20483 => "0000000000000000",20484 => "0000000000000000",
20485 => "0000000000000000",20486 => "0000000000000000",
20487 => "0000000000000000",20488 => "0000000000000000",
20489 => "0000000000000000",20490 => "0000000000000000",
20491 => "0000000000000000",20492 => "0000000000000000",
20493 => "0000000000000000",20494 => "0000000000000000",
20495 => "0000000000000000",20496 => "0000000000000000",
20497 => "0000000000000000",20498 => "0000000000000000",
20499 => "0000000000000000",20500 => "0000000000000000",
20501 => "0000000000000000",20502 => "0000000000000000",
20503 => "0000000000000000",20504 => "0000000000000000",
20505 => "0000000000000000",20506 => "0000000000000000",
20507 => "0000000000000000",20508 => "0000000000000000",
20509 => "0000000000000000",20510 => "0000000000000000",
20511 => "0000000000000000",20512 => "0000000000000000",
20513 => "0000000000000000",20514 => "0000000000000000",
20515 => "0000000000000000",20516 => "0000000000000000",
20517 => "0000000000000000",20518 => "0000000000000000",
20519 => "0000000000000000",20520 => "0000000000000000",
20521 => "0000000000000000",20522 => "0000000000000000",
20523 => "0000000000000000",20524 => "0000000000000000",
20525 => "0000000000000000",20526 => "0000000000000000",
20527 => "0000000000000000",20528 => "0000000000000000",
20529 => "0000000000000000",20530 => "0000000000000000",
20531 => "0000000000000000",20532 => "0000000000000000",
20533 => "0000000000000000",20534 => "0000000000000000",
20535 => "0000000000000000",20536 => "0000000000000000",
20537 => "0000000000000000",20538 => "0000000000000000",
20539 => "0000000000000000",20540 => "0000000000000000",
20541 => "0000000000000000",20542 => "0000000000000000",
20543 => "0000000000000000",20544 => "0000000000000000",
20545 => "0000000000000000",20546 => "0000000000000000",
20547 => "0000000000000000",20548 => "0000000000000000",
20549 => "0000000000000000",20550 => "0000000000000000",
20551 => "0000000000000000",20552 => "0000000000000000",
20553 => "0000000000000000",20554 => "0000000000000000",
20555 => "0000000000000000",20556 => "0000000000000000",
20557 => "0000000000000000",20558 => "0000000000000000",
20559 => "0000000000000000",20560 => "0000000000000000",
20561 => "0000000000000000",20562 => "0000000000000000",
20563 => "0000000000000000",20564 => "0000000000000000",
20565 => "0000000000000000",20566 => "0000000000000000",
20567 => "0000000000000000",20568 => "0000000000000000",
20569 => "0000000000000000",20570 => "0000000000000000",
20571 => "0000000000000000",20572 => "0000000000000000",
20573 => "0000000000000000",20574 => "0000000000000000",
20575 => "0000000000000000",20576 => "0000000000000000",
20577 => "0000000000000000",20578 => "0000000000000000",
20579 => "0000000000000000",20580 => "0000000000000000",
20581 => "0000000000000000",20582 => "0000000000000000",
20583 => "0000000000000000",20584 => "0000000000000000",
20585 => "0000000000000000",20586 => "0000000000000000",
20587 => "0000000000000000",20588 => "0000000000000000",
20589 => "0000000000000000",20590 => "0000000000000000",
20591 => "0000000000000000",20592 => "0000000000000000",
20593 => "0000000000000000",20594 => "0000000000000000",
20595 => "0000000000000000",20596 => "0000000000000000",
20597 => "0000000000000000",20598 => "0000000000000000",
20599 => "0000000000000000",20600 => "0000000000000000",
20601 => "0000000000000000",20602 => "0000000000000000",
20603 => "0000000000000000",20604 => "0000000000000000",
20605 => "0000000000000000",20606 => "0000000000000000",
20607 => "0000000000000000",20608 => "0000000000000000",
20609 => "0000000000000000",20610 => "0000000000000000",
20611 => "0000000000000000",20612 => "0000000000000000",
20613 => "0000000000000000",20614 => "0000000000000000",
20615 => "0000000000000000",20616 => "0000000000000000",
20617 => "0000000000000000",20618 => "0000000000000000",
20619 => "0000000000000000",20620 => "0000000000000000",
20621 => "0000000000000000",20622 => "0000000000000000",
20623 => "0000000000000000",20624 => "0000000000000000",
20625 => "0000000000000000",20626 => "0000000000000000",
20627 => "0000000000000000",20628 => "0000000000000000",
20629 => "0000000000000000",20630 => "0000000000000000",
20631 => "0000000000000000",20632 => "0000000000000000",
20633 => "0000000000000000",20634 => "0000000000000000",
20635 => "0000000000000000",20636 => "0000000000000000",
20637 => "0000000000000000",20638 => "0000000000000000",
20639 => "0000000000000000",20640 => "0000000000000000",
20641 => "0000000000000000",20642 => "0000000000000000",
20643 => "0000000000000000",20644 => "0000000000000000",
20645 => "0000000000000000",20646 => "0000000000000000",
20647 => "0000000000000000",20648 => "0000000000000000",
20649 => "0000000000000000",20650 => "0000000000000000",
20651 => "0000000000000000",20652 => "0000000000000000",
20653 => "0000000000000000",20654 => "0000000000000000",
20655 => "0000000000000000",20656 => "0000000000000000",
20657 => "0000000000000000",20658 => "0000000000000000",
20659 => "0000000000000000",20660 => "0000000000000000",
20661 => "0000000000000000",20662 => "0000000000000000",
20663 => "0000000000000000",20664 => "0000000000000000",
20665 => "0000000000000000",20666 => "0000000000000000",
20667 => "0000000000000000",20668 => "0000000000000000",
20669 => "0000000000000000",20670 => "0000000000000000",
20671 => "0000000000000000",20672 => "0000000000000000",
20673 => "0000000000000000",20674 => "0000000000000000",
20675 => "0000000000000000",20676 => "0000000000000000",
20677 => "0000000000000000",20678 => "0000000000000000",
20679 => "0000000000000000",20680 => "0000000000000000",
20681 => "0000000000000000",20682 => "0000000000000000",
20683 => "0000000000000000",20684 => "0000000000000000",
20685 => "0000000000000000",20686 => "0000000000000000",
20687 => "0000000000000000",20688 => "0000000000000000",
20689 => "0000000000000000",20690 => "0000000000000000",
20691 => "0000000000000000",20692 => "0000000000000000",
20693 => "0000000000000000",20694 => "0000000000000000",
20695 => "0000000000000000",20696 => "0000000000000000",
20697 => "0000000000000000",20698 => "0000000000000000",
20699 => "0000000000000000",20700 => "0000000000000000",
20701 => "0000000000000000",20702 => "0000000000000000",
20703 => "0000000000000000",20704 => "0000000000000000",
20705 => "0000000000000000",20706 => "0000000000000000",
20707 => "0000000000000000",20708 => "0000000000000000",
20709 => "0000000000000000",20710 => "0000000000000000",
20711 => "0000000000000000",20712 => "0000000000000000",
20713 => "0000000000000000",20714 => "0000000000000000",
20715 => "0000000000000000",20716 => "0000000000000000",
20717 => "0000000000000000",20718 => "0000000000000000",
20719 => "0000000000000000",20720 => "0000000000000000",
20721 => "0000000000000000",20722 => "0000000000000000",
20723 => "0000000000000000",20724 => "0000000000000000",
20725 => "0000000000000000",20726 => "0000000000000000",
20727 => "0000000000000000",20728 => "0000000000000000",
20729 => "0000000000000000",20730 => "0000000000000000",
20731 => "0000000000000000",20732 => "0000000000000000",
20733 => "0000000000000000",20734 => "0000000000000000",
20735 => "0000000000000000",20736 => "0000000000000000",
20737 => "0000000000000000",20738 => "0000000000000000",
20739 => "0000000000000000",20740 => "0000000000000000",
20741 => "0000000000000000",20742 => "0000000000000000",
20743 => "0000000000000000",20744 => "0000000000000000",
20745 => "0000000000000000",20746 => "0000000000000000",
20747 => "0000000000000000",20748 => "0000000000000000",
20749 => "0000000000000000",20750 => "0000000000000000",
20751 => "0000000000000000",20752 => "0000000000000000",
20753 => "0000000000000000",20754 => "0000000000000000",
20755 => "0000000000000000",20756 => "0000000000000000",
20757 => "0000000000000000",20758 => "0000000000000000",
20759 => "0000000000000000",20760 => "0000000000000000",
20761 => "0000000000000000",20762 => "0000000000000000",
20763 => "0000000000000000",20764 => "0000000000000000",
20765 => "0000000000000000",20766 => "0000000000000000",
20767 => "0000000000000000",20768 => "0000000000000000",
20769 => "0000000000000000",20770 => "0000000000000000",
20771 => "0000000000000000",20772 => "0000000000000000",
20773 => "0000000000000000",20774 => "0000000000000000",
20775 => "0000000000000000",20776 => "0000000000000000",
20777 => "0000000000000000",20778 => "0000000000000000",
20779 => "0000000000000000",20780 => "0000000000000000",
20781 => "0000000000000000",20782 => "0000000000000000",
20783 => "0000000000000000",20784 => "0000000000000000",
20785 => "0000000000000000",20786 => "0000000000000000",
20787 => "0000000000000000",20788 => "0000000000000000",
20789 => "0000000000000000",20790 => "0000000000000000",
20791 => "0000000000000000",20792 => "0000000000000000",
20793 => "0000000000000000",20794 => "0000000000000000",
20795 => "0000000000000000",20796 => "0000000000000000",
20797 => "0000000000000000",20798 => "0000000000000000",
20799 => "0000000000000000",20800 => "0000000000000000",
20801 => "0000000000000000",20802 => "0000000000000000",
20803 => "0000000000000000",20804 => "0000000000000000",
20805 => "0000000000000000",20806 => "0000000000000000",
20807 => "0000000000000000",20808 => "0000000000000000",
20809 => "0000000000000000",20810 => "0000000000000000",
20811 => "0000000000000000",20812 => "0000000000000000",
20813 => "0000000000000000",20814 => "0000000000000000",
20815 => "0000000000000000",20816 => "0000000000000000",
20817 => "0000000000000000",20818 => "0000000000000000",
20819 => "0000000000000000",20820 => "0000000000000000",
20821 => "0000000000000000",20822 => "0000000000000000",
20823 => "0000000000000000",20824 => "0000000000000000",
20825 => "0000000000000000",20826 => "0000000000000000",
20827 => "0000000000000000",20828 => "0000000000000000",
20829 => "0000000000000000",20830 => "0000000000000000",
20831 => "0000000000000000",20832 => "0000000000000000",
20833 => "0000000000000000",20834 => "0000000000000000",
20835 => "0000000000000000",20836 => "0000000000000000",
20837 => "0000000000000000",20838 => "0000000000000000",
20839 => "0000000000000000",20840 => "0000000000000000",
20841 => "0000000000000000",20842 => "0000000000000000",
20843 => "0000000000000000",20844 => "0000000000000000",
20845 => "0000000000000000",20846 => "0000000000000000",
20847 => "0000000000000000",20848 => "0000000000000000",
20849 => "0000000000000000",20850 => "0000000000000000",
20851 => "0000000000000000",20852 => "0000000000000000",
20853 => "0000000000000000",20854 => "0000000000000000",
20855 => "0000000000000000",20856 => "0000000000000000",
20857 => "0000000000000000",20858 => "0000000000000000",
20859 => "0000000000000000",20860 => "0000000000000000",
20861 => "0000000000000000",20862 => "0000000000000000",
20863 => "0000000000000000",20864 => "0000000000000000",
20865 => "0000000000000000",20866 => "0000000000000000",
20867 => "0000000000000000",20868 => "0000000000000000",
20869 => "0000000000000000",20870 => "0000000000000000",
20871 => "0000000000000000",20872 => "0000000000000000",
20873 => "0000000000000000",20874 => "0000000000000000",
20875 => "0000000000000000",20876 => "0000000000000000",
20877 => "0000000000000000",20878 => "0000000000000000",
20879 => "0000000000000000",20880 => "0000000000000000",
20881 => "0000000000000000",20882 => "0000000000000000",
20883 => "0000000000000000",20884 => "0000000000000000",
20885 => "0000000000000000",20886 => "0000000000000000",
20887 => "0000000000000000",20888 => "0000000000000000",
20889 => "0000000000000000",20890 => "0000000000000000",
20891 => "0000000000000000",20892 => "0000000000000000",
20893 => "0000000000000000",20894 => "0000000000000000",
20895 => "0000000000000000",20896 => "0000000000000000",
20897 => "0000000000000000",20898 => "0000000000000000",
20899 => "0000000000000000",20900 => "0000000000000000",
20901 => "0000000000000000",20902 => "0000000000000000",
20903 => "0000000000000000",20904 => "0000000000000000",
20905 => "0000000000000000",20906 => "0000000000000000",
20907 => "0000000000000000",20908 => "0000000000000000",
20909 => "0000000000000000",20910 => "0000000000000000",
20911 => "0000000000000000",20912 => "0000000000000000",
20913 => "0000000000000000",20914 => "0000000000000000",
20915 => "0000000000000000",20916 => "0000000000000000",
20917 => "0000000000000000",20918 => "0000000000000000",
20919 => "0000000000000000",20920 => "0000000000000000",
20921 => "0000000000000000",20922 => "0000000000000000",
20923 => "0000000000000000",20924 => "0000000000000000",
20925 => "0000000000000000",20926 => "0000000000000000",
20927 => "0000000000000000",20928 => "0000000000000000",
20929 => "0000000000000000",20930 => "0000000000000000",
20931 => "0000000000000000",20932 => "0000000000000000",
20933 => "0000000000000000",20934 => "0000000000000000",
20935 => "0000000000000000",20936 => "0000000000000000",
20937 => "0000000000000000",20938 => "0000000000000000",
20939 => "0000000000000000",20940 => "0000000000000000",
20941 => "0000000000000000",20942 => "0000000000000000",
20943 => "0000000000000000",20944 => "0000000000000000",
20945 => "0000000000000000",20946 => "0000000000000000",
20947 => "0000000000000000",20948 => "0000000000000000",
20949 => "0000000000000000",20950 => "0000000000000000",
20951 => "0000000000000000",20952 => "0000000000000000",
20953 => "0000000000000000",20954 => "0000000000000000",
20955 => "0000000000000000",20956 => "0000000000000000",
20957 => "0000000000000000",20958 => "0000000000000000",
20959 => "0000000000000000",20960 => "0000000000000000",
20961 => "0000000000000000",20962 => "0000000000000000",
20963 => "0000000000000000",20964 => "0000000000000000",
20965 => "0000000000000000",20966 => "0000000000000000",
20967 => "0000000000000000",20968 => "0000000000000000",
20969 => "0000000000000000",20970 => "0000000000000000",
20971 => "0000000000000000",20972 => "0000000000000000",
20973 => "0000000000000000",20974 => "0000000000000000",
20975 => "0000000000000000",20976 => "0000000000000000",
20977 => "0000000000000000",20978 => "0000000000000000",
20979 => "0000000000000000",20980 => "0000000000000000",
20981 => "0000000000000000",20982 => "0000000000000000",
20983 => "0000000000000000",20984 => "0000000000000000",
20985 => "0000000000000000",20986 => "0000000000000000",
20987 => "0000000000000000",20988 => "0000000000000000",
20989 => "0000000000000000",20990 => "0000000000000000",
20991 => "0000000000000000",20992 => "0000000000000000",
20993 => "0000000000000000",20994 => "0000000000000000",
20995 => "0000000000000000",20996 => "0000000000000000",
20997 => "0000000000000000",20998 => "0000000000000000",
20999 => "0000000000000000",21000 => "0000000000000000",
21001 => "0000000000000000",21002 => "0000000000000000",
21003 => "0000000000000000",21004 => "0000000000000000",
21005 => "0000000000000000",21006 => "0000000000000000",
21007 => "0000000000000000",21008 => "0000000000000000",
21009 => "0000000000000000",21010 => "0000000000000000",
21011 => "0000000000000000",21012 => "0000000000000000",
21013 => "0000000000000000",21014 => "0000000000000000",
21015 => "0000000000000000",21016 => "0000000000000000",
21017 => "0000000000000000",21018 => "0000000000000000",
21019 => "0000000000000000",21020 => "0000000000000000",
21021 => "0000000000000000",21022 => "0000000000000000",
21023 => "0000000000000000",21024 => "0000000000000000",
21025 => "0000000000000000",21026 => "0000000000000000",
21027 => "0000000000000000",21028 => "0000000000000000",
21029 => "0000000000000000",21030 => "0000000000000000",
21031 => "0000000000000000",21032 => "0000000000000000",
21033 => "0000000000000000",21034 => "0000000000000000",
21035 => "0000000000000000",21036 => "0000000000000000",
21037 => "0000000000000000",21038 => "0000000000000000",
21039 => "0000000000000000",21040 => "0000000000000000",
21041 => "0000000000000000",21042 => "0000000000000000",
21043 => "0000000000000000",21044 => "0000000000000000",
21045 => "0000000000000000",21046 => "0000000000000000",
21047 => "0000000000000000",21048 => "0000000000000000",
21049 => "0000000000000000",21050 => "0000000000000000",
21051 => "0000000000000000",21052 => "0000000000000000",
21053 => "0000000000000000",21054 => "0000000000000000",
21055 => "0000000000000000",21056 => "0000000000000000",
21057 => "0000000000000000",21058 => "0000000000000000",
21059 => "0000000000000000",21060 => "0000000000000000",
21061 => "0000000000000000",21062 => "0000000000000000",
21063 => "0000000000000000",21064 => "0000000000000000",
21065 => "0000000000000000",21066 => "0000000000000000",
21067 => "0000000000000000",21068 => "0000000000000000",
21069 => "0000000000000000",21070 => "0000000000000000",
21071 => "0000000000000000",21072 => "0000000000000000",
21073 => "0000000000000000",21074 => "0000000000000000",
21075 => "0000000000000000",21076 => "0000000000000000",
21077 => "0000000000000000",21078 => "0000000000000000",
21079 => "0000000000000000",21080 => "0000000000000000",
21081 => "0000000000000000",21082 => "0000000000000000",
21083 => "0000000000000000",21084 => "0000000000000000",
21085 => "0000000000000000",21086 => "0000000000000000",
21087 => "0000000000000000",21088 => "0000000000000000",
21089 => "0000000000000000",21090 => "0000000000000000",
21091 => "0000000000000000",21092 => "0000000000000000",
21093 => "0000000000000000",21094 => "0000000000000000",
21095 => "0000000000000000",21096 => "0000000000000000",
21097 => "0000000000000000",21098 => "0000000000000000",
21099 => "0000000000000000",21100 => "0000000000000000",
21101 => "0000000000000000",21102 => "0000000000000000",
21103 => "0000000000000000",21104 => "0000000000000000",
21105 => "0000000000000000",21106 => "0000000000000000",
21107 => "0000000000000000",21108 => "0000000000000000",
21109 => "0000000000000000",21110 => "0000000000000000",
21111 => "0000000000000000",21112 => "0000000000000000",
21113 => "0000000000000000",21114 => "0000000000000000",
21115 => "0000000000000000",21116 => "0000000000000000",
21117 => "0000000000000000",21118 => "0000000000000000",
21119 => "0000000000000000",21120 => "0000000000000000",
21121 => "0000000000000000",21122 => "0000000000000000",
21123 => "0000000000000000",21124 => "0000000000000000",
21125 => "0000000000000000",21126 => "0000000000000000",
21127 => "0000000000000000",21128 => "0000000000000000",
21129 => "0000000000000000",21130 => "0000000000000000",
21131 => "0000000000000000",21132 => "0000000000000000",
21133 => "0000000000000000",21134 => "0000000000000000",
21135 => "0000000000000000",21136 => "0000000000000000",
21137 => "0000000000000000",21138 => "0000000000000000",
21139 => "0000000000000000",21140 => "0000000000000000",
21141 => "0000000000000000",21142 => "0000000000000000",
21143 => "0000000000000000",21144 => "0000000000000000",
21145 => "0000000000000000",21146 => "0000000000000000",
21147 => "0000000000000000",21148 => "0000000000000000",
21149 => "0000000000000000",21150 => "0000000000000000",
21151 => "0000000000000000",21152 => "0000000000000000",
21153 => "0000000000000000",21154 => "0000000000000000",
21155 => "0000000000000000",21156 => "0000000000000000",
21157 => "0000000000000000",21158 => "0000000000000000",
21159 => "0000000000000000",21160 => "0000000000000000",
21161 => "0000000000000000",21162 => "0000000000000000",
21163 => "0000000000000000",21164 => "0000000000000000",
21165 => "0000000000000000",21166 => "0000000000000000",
21167 => "0000000000000000",21168 => "0000000000000000",
21169 => "0000000000000000",21170 => "0000000000000000",
21171 => "0000000000000000",21172 => "0000000000000000",
21173 => "0000000000000000",21174 => "0000000000000000",
21175 => "0000000000000000",21176 => "0000000000000000",
21177 => "0000000000000000",21178 => "0000000000000000",
21179 => "0000000000000000",21180 => "0000000000000000",
21181 => "0000000000000000",21182 => "0000000000000000",
21183 => "0000000000000000",21184 => "0000000000000000",
21185 => "0000000000000000",21186 => "0000000000000000",
21187 => "0000000000000000",21188 => "0000000000000000",
21189 => "0000000000000000",21190 => "0000000000000000",
21191 => "0000000000000000",21192 => "0000000000000000",
21193 => "0000000000000000",21194 => "0000000000000000",
21195 => "0000000000000000",21196 => "0000000000000000",
21197 => "0000000000000000",21198 => "0000000000000000",
21199 => "0000000000000000",21200 => "0000000000000000",
21201 => "0000000000000000",21202 => "0000000000000000",
21203 => "0000000000000000",21204 => "0000000000000000",
21205 => "0000000000000000",21206 => "0000000000000000",
21207 => "0000000000000000",21208 => "0000000000000000",
21209 => "0000000000000000",21210 => "0000000000000000",
21211 => "0000000000000000",21212 => "0000000000000000",
21213 => "0000000000000000",21214 => "0000000000000000",
21215 => "0000000000000000",21216 => "0000000000000000",
21217 => "0000000000000000",21218 => "0000000000000000",
21219 => "0000000000000000",21220 => "0000000000000000",
21221 => "0000000000000000",21222 => "0000000000000000",
21223 => "0000000000000000",21224 => "0000000000000000",
21225 => "0000000000000000",21226 => "0000000000000000",
21227 => "0000000000000000",21228 => "0000000000000000",
21229 => "0000000000000000",21230 => "0000000000000000",
21231 => "0000000000000000",21232 => "0000000000000000",
21233 => "0000000000000000",21234 => "0000000000000000",
21235 => "0000000000000000",21236 => "0000000000000000",
21237 => "0000000000000000",21238 => "0000000000000000",
21239 => "0000000000000000",21240 => "0000000000000000",
21241 => "0000000000000000",21242 => "0000000000000000",
21243 => "0000000000000000",21244 => "0000000000000000",
21245 => "0000000000000000",21246 => "0000000000000000",
21247 => "0000000000000000",21248 => "0000000000000000",
21249 => "0000000000000000",21250 => "0000000000000000",
21251 => "0000000000000000",21252 => "0000000000000000",
21253 => "0000000000000000",21254 => "0000000000000000",
21255 => "0000000000000000",21256 => "0000000000000000",
21257 => "0000000000000000",21258 => "0000000000000000",
21259 => "0000000000000000",21260 => "0000000000000000",
21261 => "0000000000000000",21262 => "0000000000000000",
21263 => "0000000000000000",21264 => "0000000000000000",
21265 => "0000000000000000",21266 => "0000000000000000",
21267 => "0000000000000000",21268 => "0000000000000000",
21269 => "0000000000000000",21270 => "0000000000000000",
21271 => "0000000000000000",21272 => "0000000000000000",
21273 => "0000000000000000",21274 => "0000000000000000",
21275 => "0000000000000000",21276 => "0000000000000000",
21277 => "0000000000000000",21278 => "0000000000000000",
21279 => "0000000000000000",21280 => "0000000000000000",
21281 => "0000000000000000",21282 => "0000000000000000",
21283 => "0000000000000000",21284 => "0000000000000000",
21285 => "0000000000000000",21286 => "0000000000000000",
21287 => "0000000000000000",21288 => "0000000000000000",
21289 => "0000000000000000",21290 => "0000000000000000",
21291 => "0000000000000000",21292 => "0000000000000000",
21293 => "0000000000000000",21294 => "0000000000000000",
21295 => "0000000000000000",21296 => "0000000000000000",
21297 => "0000000000000000",21298 => "0000000000000000",
21299 => "0000000000000000",21300 => "0000000000000000",
21301 => "0000000000000000",21302 => "0000000000000000",
21303 => "0000000000000000",21304 => "0000000000000000",
21305 => "0000000000000000",21306 => "0000000000000000",
21307 => "0000000000000000",21308 => "0000000000000000",
21309 => "0000000000000000",21310 => "0000000000000000",
21311 => "0000000000000000",21312 => "0000000000000000",
21313 => "0000000000000000",21314 => "0000000000000000",
21315 => "0000000000000000",21316 => "0000000000000000",
21317 => "0000000000000000",21318 => "0000000000000000",
21319 => "0000000000000000",21320 => "0000000000000000",
21321 => "0000000000000000",21322 => "0000000000000000",
21323 => "0000000000000000",21324 => "0000000000000000",
21325 => "0000000000000000",21326 => "0000000000000000",
21327 => "0000000000000000",21328 => "0000000000000000",
21329 => "0000000000000000",21330 => "0000000000000000",
21331 => "0000000000000000",21332 => "0000000000000000",
21333 => "0000000000000000",21334 => "0000000000000000",
21335 => "0000000000000000",21336 => "0000000000000000",
21337 => "0000000000000000",21338 => "0000000000000000",
21339 => "0000000000000000",21340 => "0000000000000000",
21341 => "0000000000000000",21342 => "0000000000000000",
21343 => "0000000000000000",21344 => "0000000000000000",
21345 => "0000000000000000",21346 => "0000000000000000",
21347 => "0000000000000000",21348 => "0000000000000000",
21349 => "0000000000000000",21350 => "0000000000000000",
21351 => "0000000000000000",21352 => "0000000000000000",
21353 => "0000000000000000",21354 => "0000000000000000",
21355 => "0000000000000000",21356 => "0000000000000000",
21357 => "0000000000000000",21358 => "0000000000000000",
21359 => "0000000000000000",21360 => "0000000000000000",
21361 => "0000000000000000",21362 => "0000000000000000",
21363 => "0000000000000000",21364 => "0000000000000000",
21365 => "0000000000000000",21366 => "0000000000000000",
21367 => "0000000000000000",21368 => "0000000000000000",
21369 => "0000000000000000",21370 => "0000000000000000",
21371 => "0000000000000000",21372 => "0000000000000000",
21373 => "0000000000000000",21374 => "0000000000000000",
21375 => "0000000000000000",21376 => "0000000000000000",
21377 => "0000000000000000",21378 => "0000000000000000",
21379 => "0000000000000000",21380 => "0000000000000000",
21381 => "0000000000000000",21382 => "0000000000000000",
21383 => "0000000000000000",21384 => "0000000000000000",
21385 => "0000000000000000",21386 => "0000000000000000",
21387 => "0000000000000000",21388 => "0000000000000000",
21389 => "0000000000000000",21390 => "0000000000000000",
21391 => "0000000000000000",21392 => "0000000000000000",
21393 => "0000000000000000",21394 => "0000000000000000",
21395 => "0000000000000000",21396 => "0000000000000000",
21397 => "0000000000000000",21398 => "0000000000000000",
21399 => "0000000000000000",21400 => "0000000000000000",
21401 => "0000000000000000",21402 => "0000000000000000",
21403 => "0000000000000000",21404 => "0000000000000000",
21405 => "0000000000000000",21406 => "0000000000000000",
21407 => "0000000000000000",21408 => "0000000000000000",
21409 => "0000000000000000",21410 => "0000000000000000",
21411 => "0000000000000000",21412 => "0000000000000000",
21413 => "0000000000000000",21414 => "0000000000000000",
21415 => "0000000000000000",21416 => "0000000000000000",
21417 => "0000000000000000",21418 => "0000000000000000",
21419 => "0000000000000000",21420 => "0000000000000000",
21421 => "0000000000000000",21422 => "0000000000000000",
21423 => "0000000000000000",21424 => "0000000000000000",
21425 => "0000000000000000",21426 => "0000000000000000",
21427 => "0000000000000000",21428 => "0000000000000000",
21429 => "0000000000000000",21430 => "0000000000000000",
21431 => "0000000000000000",21432 => "0000000000000000",
21433 => "0000000000000000",21434 => "0000000000000000",
21435 => "0000000000000000",21436 => "0000000000000000",
21437 => "0000000000000000",21438 => "0000000000000000",
21439 => "0000000000000000",21440 => "0000000000000000",
21441 => "0000000000000000",21442 => "0000000000000000",
21443 => "0000000000000000",21444 => "0000000000000000",
21445 => "0000000000000000",21446 => "0000000000000000",
21447 => "0000000000000000",21448 => "0000000000000000",
21449 => "0000000000000000",21450 => "0000000000000000",
21451 => "0000000000000000",21452 => "0000000000000000",
21453 => "0000000000000000",21454 => "0000000000000000",
21455 => "0000000000000000",21456 => "0000000000000000",
21457 => "0000000000000000",21458 => "0000000000000000",
21459 => "0000000000000000",21460 => "0000000000000000",
21461 => "0000000000000000",21462 => "0000000000000000",
21463 => "0000000000000000",21464 => "0000000000000000",
21465 => "0000000000000000",21466 => "0000000000000000",
21467 => "0000000000000000",21468 => "0000000000000000",
21469 => "0000000000000000",21470 => "0000000000000000",
21471 => "0000000000000000",21472 => "0000000000000000",
21473 => "0000000000000000",21474 => "0000000000000000",
21475 => "0000000000000000",21476 => "0000000000000000",
21477 => "0000000000000000",21478 => "0000000000000000",
21479 => "0000000000000000",21480 => "0000000000000000",
21481 => "0000000000000000",21482 => "0000000000000000",
21483 => "0000000000000000",21484 => "0000000000000000",
21485 => "0000000000000000",21486 => "0000000000000000",
21487 => "0000000000000000",21488 => "0000000000000000",
21489 => "0000000000000000",21490 => "0000000000000000",
21491 => "0000000000000000",21492 => "0000000000000000",
21493 => "0000000000000000",21494 => "0000000000000000",
21495 => "0000000000000000",21496 => "0000000000000000",
21497 => "0000000000000000",21498 => "0000000000000000",
21499 => "0000000000000000",21500 => "0000000000000000",
21501 => "0000000000000000",21502 => "0000000000000000",
21503 => "0000000000000000",21504 => "0000000000000000",
21505 => "0000000000000000",21506 => "0000000000000000",
21507 => "0000000000000000",21508 => "0000000000000000",
21509 => "0000000000000000",21510 => "0000000000000000",
21511 => "0000000000000000",21512 => "0000000000000000",
21513 => "0000000000000000",21514 => "0000000000000000",
21515 => "0000000000000000",21516 => "0000000000000000",
21517 => "0000000000000000",21518 => "0000000000000000",
21519 => "0000000000000000",21520 => "0000000000000000",
21521 => "0000000000000000",21522 => "0000000000000000",
21523 => "0000000000000000",21524 => "0000000000000000",
21525 => "0000000000000000",21526 => "0000000000000000",
21527 => "0000000000000000",21528 => "0000000000000000",
21529 => "0000000000000000",21530 => "0000000000000000",
21531 => "0000000000000000",21532 => "0000000000000000",
21533 => "0000000000000000",21534 => "0000000000000000",
21535 => "0000000000000000",21536 => "0000000000000000",
21537 => "0000000000000000",21538 => "0000000000000000",
21539 => "0000000000000000",21540 => "0000000000000000",
21541 => "0000000000000000",21542 => "0000000000000000",
21543 => "0000000000000000",21544 => "0000000000000000",
21545 => "0000000000000000",21546 => "0000000000000000",
21547 => "0000000000000000",21548 => "0000000000000000",
21549 => "0000000000000000",21550 => "0000000000000000",
21551 => "0000000000000000",21552 => "0000000000000000",
21553 => "0000000000000000",21554 => "0000000000000000",
21555 => "0000000000000000",21556 => "0000000000000000",
21557 => "0000000000000000",21558 => "0000000000000000",
21559 => "0000000000000000",21560 => "0000000000000000",
21561 => "0000000000000000",21562 => "0000000000000000",
21563 => "0000000000000000",21564 => "0000000000000000",
21565 => "0000000000000000",21566 => "0000000000000000",
21567 => "0000000000000000",21568 => "0000000000000000",
21569 => "0000000000000000",21570 => "0000000000000000",
21571 => "0000000000000000",21572 => "0000000000000000",
21573 => "0000000000000000",21574 => "0000000000000000",
21575 => "0000000000000000",21576 => "0000000000000000",
21577 => "0000000000000000",21578 => "0000000000000000",
21579 => "0000000000000000",21580 => "0000000000000000",
21581 => "0000000000000000",21582 => "0000000000000000",
21583 => "0000000000000000",21584 => "0000000000000000",
21585 => "0000000000000000",21586 => "0000000000000000",
21587 => "0000000000000000",21588 => "0000000000000000",
21589 => "0000000000000000",21590 => "0000000000000000",
21591 => "0000000000000000",21592 => "0000000000000000",
21593 => "0000000000000000",21594 => "0000000000000000",
21595 => "0000000000000000",21596 => "0000000000000000",
21597 => "0000000000000000",21598 => "0000000000000000",
21599 => "0000000000000000",21600 => "0000000000000000",
21601 => "0000000000000000",21602 => "0000000000000000",
21603 => "0000000000000000",21604 => "0000000000000000",
21605 => "0000000000000000",21606 => "0000000000000000",
21607 => "0000000000000000",21608 => "0000000000000000",
21609 => "0000000000000000",21610 => "0000000000000000",
21611 => "0000000000000000",21612 => "0000000000000000",
21613 => "0000000000000000",21614 => "0000000000000000",
21615 => "0000000000000000",21616 => "0000000000000000",
21617 => "0000000000000000",21618 => "0000000000000000",
21619 => "0000000000000000",21620 => "0000000000000000",
21621 => "0000000000000000",21622 => "0000000000000000",
21623 => "0000000000000000",21624 => "0000000000000000",
21625 => "0000000000000000",21626 => "0000000000000000",
21627 => "0000000000000000",21628 => "0000000000000000",
21629 => "0000000000000000",21630 => "0000000000000000",
21631 => "0000000000000000",21632 => "0000000000000000",
21633 => "0000000000000000",21634 => "0000000000000000",
21635 => "0000000000000000",21636 => "0000000000000000",
21637 => "0000000000000000",21638 => "0000000000000000",
21639 => "0000000000000000",21640 => "0000000000000000",
21641 => "0000000000000000",21642 => "0000000000000000",
21643 => "0000000000000000",21644 => "0000000000000000",
21645 => "0000000000000000",21646 => "0000000000000000",
21647 => "0000000000000000",21648 => "0000000000000000",
21649 => "0000000000000000",21650 => "0000000000000000",
21651 => "0000000000000000",21652 => "0000000000000000",
21653 => "0000000000000000",21654 => "0000000000000000",
21655 => "0000000000000000",21656 => "0000000000000000",
21657 => "0000000000000000",21658 => "0000000000000000",
21659 => "0000000000000000",21660 => "0000000000000000",
21661 => "0000000000000000",21662 => "0000000000000000",
21663 => "0000000000000000",21664 => "0000000000000000",
21665 => "0000000000000000",21666 => "0000000000000000",
21667 => "0000000000000000",21668 => "0000000000000000",
21669 => "0000000000000000",21670 => "0000000000000000",
21671 => "0000000000000000",21672 => "0000000000000000",
21673 => "0000000000000000",21674 => "0000000000000000",
21675 => "0000000000000000",21676 => "0000000000000000",
21677 => "0000000000000000",21678 => "0000000000000000",
21679 => "0000000000000000",21680 => "0000000000000000",
21681 => "0000000000000000",21682 => "0000000000000000",
21683 => "0000000000000000",21684 => "0000000000000000",
21685 => "0000000000000000",21686 => "0000000000000000",
21687 => "0000000000000000",21688 => "0000000000000000",
21689 => "0000000000000000",21690 => "0000000000000000",
21691 => "0000000000000000",21692 => "0000000000000000",
21693 => "0000000000000000",21694 => "0000000000000000",
21695 => "0000000000000000",21696 => "0000000000000000",
21697 => "0000000000000000",21698 => "0000000000000000",
21699 => "0000000000000000",21700 => "0000000000000000",
21701 => "0000000000000000",21702 => "0000000000000000",
21703 => "0000000000000000",21704 => "0000000000000000",
21705 => "0000000000000000",21706 => "0000000000000000",
21707 => "0000000000000000",21708 => "0000000000000000",
21709 => "0000000000000000",21710 => "0000000000000000",
21711 => "0000000000000000",21712 => "0000000000000000",
21713 => "0000000000000000",21714 => "0000000000000000",
21715 => "0000000000000000",21716 => "0000000000000000",
21717 => "0000000000000000",21718 => "0000000000000000",
21719 => "0000000000000000",21720 => "0000000000000000",
21721 => "0000000000000000",21722 => "0000000000000000",
21723 => "0000000000000000",21724 => "0000000000000000",
21725 => "0000000000000000",21726 => "0000000000000000",
21727 => "0000000000000000",21728 => "0000000000000000",
21729 => "0000000000000000",21730 => "0000000000000000",
21731 => "0000000000000000",21732 => "0000000000000000",
21733 => "0000000000000000",21734 => "0000000000000000",
21735 => "0000000000000000",21736 => "0000000000000000",
21737 => "0000000000000000",21738 => "0000000000000000",
21739 => "0000000000000000",21740 => "0000000000000000",
21741 => "0000000000000000",21742 => "0000000000000000",
21743 => "0000000000000000",21744 => "0000000000000000",
21745 => "0000000000000000",21746 => "0000000000000000",
21747 => "0000000000000000",21748 => "0000000000000000",
21749 => "0000000000000000",21750 => "0000000000000000",
21751 => "0000000000000000",21752 => "0000000000000000",
21753 => "0000000000000000",21754 => "0000000000000000",
21755 => "0000000000000000",21756 => "0000000000000000",
21757 => "0000000000000000",21758 => "0000000000000000",
21759 => "0000000000000000",21760 => "0000000000000000",
21761 => "0000000000000000",21762 => "0000000000000000",
21763 => "0000000000000000",21764 => "0000000000000000",
21765 => "0000000000000000",21766 => "0000000000000000",
21767 => "0000000000000000",21768 => "0000000000000000",
21769 => "0000000000000000",21770 => "0000000000000000",
21771 => "0000000000000000",21772 => "0000000000000000",
21773 => "0000000000000000",21774 => "0000000000000000",
21775 => "0000000000000000",21776 => "0000000000000000",
21777 => "0000000000000000",21778 => "0000000000000000",
21779 => "0000000000000000",21780 => "0000000000000000",
21781 => "0000000000000000",21782 => "0000000000000000",
21783 => "0000000000000000",21784 => "0000000000000000",
21785 => "0000000000000000",21786 => "0000000000000000",
21787 => "0000000000000000",21788 => "0000000000000000",
21789 => "0000000000000000",21790 => "0000000000000000",
21791 => "0000000000000000",21792 => "0000000000000000",
21793 => "0000000000000000",21794 => "0000000000000000",
21795 => "0000000000000000",21796 => "0000000000000000",
21797 => "0000000000000000",21798 => "0000000000000000",
21799 => "0000000000000000",21800 => "0000000000000000",
21801 => "0000000000000000",21802 => "0000000000000000",
21803 => "0000000000000000",21804 => "0000000000000000",
21805 => "0000000000000000",21806 => "0000000000000000",
21807 => "0000000000000000",21808 => "0000000000000000",
21809 => "0000000000000000",21810 => "0000000000000000",
21811 => "0000000000000000",21812 => "0000000000000000",
21813 => "0000000000000000",21814 => "0000000000000000",
21815 => "0000000000000000",21816 => "0000000000000000",
21817 => "0000000000000000",21818 => "0000000000000000",
21819 => "0000000000000000",21820 => "0000000000000000",
21821 => "0000000000000000",21822 => "0000000000000000",
21823 => "0000000000000000",21824 => "0000000000000000",
21825 => "0000000000000000",21826 => "0000000000000000",
21827 => "0000000000000000",21828 => "0000000000000000",
21829 => "0000000000000000",21830 => "0000000000000000",
21831 => "0000000000000000",21832 => "0000000000000000",
21833 => "0000000000000000",21834 => "0000000000000000",
21835 => "0000000000000000",21836 => "0000000000000000",
21837 => "0000000000000000",21838 => "0000000000000000",
21839 => "0000000000000000",21840 => "0000000000000000",
21841 => "0000000000000000",21842 => "0000000000000000",
21843 => "0000000000000000",21844 => "0000000000000000",
21845 => "0000000000000000",21846 => "0000000000000000",
21847 => "0000000000000000",21848 => "0000000000000000",
21849 => "0000000000000000",21850 => "0000000000000000",
21851 => "0000000000000000",21852 => "0000000000000000",
21853 => "0000000000000000",21854 => "0000000000000000",
21855 => "0000000000000000",21856 => "0000000000000000",
21857 => "0000000000000000",21858 => "0000000000000000",
21859 => "0000000000000000",21860 => "0000000000000000",
21861 => "0000000000000000",21862 => "0000000000000000",
21863 => "0000000000000000",21864 => "0000000000000000",
21865 => "0000000000000000",21866 => "0000000000000000",
21867 => "0000000000000000",21868 => "0000000000000000",
21869 => "0000000000000000",21870 => "0000000000000000",
21871 => "0000000000000000",21872 => "0000000000000000",
21873 => "0000000000000000",21874 => "0000000000000000",
21875 => "0000000000000000",21876 => "0000000000000000",
21877 => "0000000000000000",21878 => "0000000000000000",
21879 => "0000000000000000",21880 => "0000000000000000",
21881 => "0000000000000000",21882 => "0000000000000000",
21883 => "0000000000000000",21884 => "0000000000000000",
21885 => "0000000000000000",21886 => "0000000000000000",
21887 => "0000000000000000",21888 => "0000000000000000",
21889 => "0000000000000000",21890 => "0000000000000000",
21891 => "0000000000000000",21892 => "0000000000000000",
21893 => "0000000000000000",21894 => "0000000000000000",
21895 => "0000000000000000",21896 => "0000000000000000",
21897 => "0000000000000000",21898 => "0000000000000000",
21899 => "0000000000000000",21900 => "0000000000000000",
21901 => "0000000000000000",21902 => "0000000000000000",
21903 => "0000000000000000",21904 => "0000000000000000",
21905 => "0000000000000000",21906 => "0000000000000000",
21907 => "0000000000000000",21908 => "0000000000000000",
21909 => "0000000000000000",21910 => "0000000000000000",
21911 => "0000000000000000",21912 => "0000000000000000",
21913 => "0000000000000000",21914 => "0000000000000000",
21915 => "0000000000000000",21916 => "0000000000000000",
21917 => "0000000000000000",21918 => "0000000000000000",
21919 => "0000000000000000",21920 => "0000000000000000",
21921 => "0000000000000000",21922 => "0000000000000000",
21923 => "0000000000000000",21924 => "0000000000000000",
21925 => "0000000000000000",21926 => "0000000000000000",
21927 => "0000000000000000",21928 => "0000000000000000",
21929 => "0000000000000000",21930 => "0000000000000000",
21931 => "0000000000000000",21932 => "0000000000000000",
21933 => "0000000000000000",21934 => "0000000000000000",
21935 => "0000000000000000",21936 => "0000000000000000",
21937 => "0000000000000000",21938 => "0000000000000000",
21939 => "0000000000000000",21940 => "0000000000000000",
21941 => "0000000000000000",21942 => "0000000000000000",
21943 => "0000000000000000",21944 => "0000000000000000",
21945 => "0000000000000000",21946 => "0000000000000000",
21947 => "0000000000000000",21948 => "0000000000000000",
21949 => "0000000000000000",21950 => "0000000000000000",
21951 => "0000000000000000",21952 => "0000000000000000",
21953 => "0000000000000000",21954 => "0000000000000000",
21955 => "0000000000000000",21956 => "0000000000000000",
21957 => "0000000000000000",21958 => "0000000000000000",
21959 => "0000000000000000",21960 => "0000000000000000",
21961 => "0000000000000000",21962 => "0000000000000000",
21963 => "0000000000000000",21964 => "0000000000000000",
21965 => "0000000000000000",21966 => "0000000000000000",
21967 => "0000000000000000",21968 => "0000000000000000",
21969 => "0000000000000000",21970 => "0000000000000000",
21971 => "0000000000000000",21972 => "0000000000000000",
21973 => "0000000000000000",21974 => "0000000000000000",
21975 => "0000000000000000",21976 => "0000000000000000",
21977 => "0000000000000000",21978 => "0000000000000000",
21979 => "0000000000000000",21980 => "0000000000000000",
21981 => "0000000000000000",21982 => "0000000000000000",
21983 => "0000000000000000",21984 => "0000000000000000",
21985 => "0000000000000000",21986 => "0000000000000000",
21987 => "0000000000000000",21988 => "0000000000000000",
21989 => "0000000000000000",21990 => "0000000000000000",
21991 => "0000000000000000",21992 => "0000000000000000",
21993 => "0000000000000000",21994 => "0000000000000000",
21995 => "0000000000000000",21996 => "0000000000000000",
21997 => "0000000000000000",21998 => "0000000000000000",
21999 => "0000000000000000",22000 => "0000000000000000",
22001 => "0000000000000000",22002 => "0000000000000000",
22003 => "0000000000000000",22004 => "0000000000000000",
22005 => "0000000000000000",22006 => "0000000000000000",
22007 => "0000000000000000",22008 => "0000000000000000",
22009 => "0000000000000000",22010 => "0000000000000000",
22011 => "0000000000000000",22012 => "0000000000000000",
22013 => "0000000000000000",22014 => "0000000000000000",
22015 => "0000000000000000",22016 => "0000000000000000",
22017 => "0000000000000000",22018 => "0000000000000000",
22019 => "0000000000000000",22020 => "0000000000000000",
22021 => "0000000000000000",22022 => "0000000000000000",
22023 => "0000000000000000",22024 => "0000000000000000",
22025 => "0000000000000000",22026 => "0000000000000000",
22027 => "0000000000000000",22028 => "0000000000000000",
22029 => "0000000000000000",22030 => "0000000000000000",
22031 => "0000000000000000",22032 => "0000000000000000",
22033 => "0000000000000000",22034 => "0000000000000000",
22035 => "0000000000000000",22036 => "0000000000000000",
22037 => "0000000000000000",22038 => "0000000000000000",
22039 => "0000000000000000",22040 => "0000000000000000",
22041 => "0000000000000000",22042 => "0000000000000000",
22043 => "0000000000000000",22044 => "0000000000000000",
22045 => "0000000000000000",22046 => "0000000000000000",
22047 => "0000000000000000",22048 => "0000000000000000",
22049 => "0000000000000000",22050 => "0000000000000000",
22051 => "0000000000000000",22052 => "0000000000000000",
22053 => "0000000000000000",22054 => "0000000000000000",
22055 => "0000000000000000",22056 => "0000000000000000",
22057 => "0000000000000000",22058 => "0000000000000000",
22059 => "0000000000000000",22060 => "0000000000000000",
22061 => "0000000000000000",22062 => "0000000000000000",
22063 => "0000000000000000",22064 => "0000000000000000",
22065 => "0000000000000000",22066 => "0000000000000000",
22067 => "0000000000000000",22068 => "0000000000000000",
22069 => "0000000000000000",22070 => "0000000000000000",
22071 => "0000000000000000",22072 => "0000000000000000",
22073 => "0000000000000000",22074 => "0000000000000000",
22075 => "0000000000000000",22076 => "0000000000000000",
22077 => "0000000000000000",22078 => "0000000000000000",
22079 => "0000000000000000",22080 => "0000000000000000",
22081 => "0000000000000000",22082 => "0000000000000000",
22083 => "0000000000000000",22084 => "0000000000000000",
22085 => "0000000000000000",22086 => "0000000000000000",
22087 => "0000000000000000",22088 => "0000000000000000",
22089 => "0000000000000000",22090 => "0000000000000000",
22091 => "0000000000000000",22092 => "0000000000000000",
22093 => "0000000000000000",22094 => "0000000000000000",
22095 => "0000000000000000",22096 => "0000000000000000",
22097 => "0000000000000000",22098 => "0000000000000000",
22099 => "0000000000000000",22100 => "0000000000000000",
22101 => "0000000000000000",22102 => "0000000000000000",
22103 => "0000000000000000",22104 => "0000000000000000",
22105 => "0000000000000000",22106 => "0000000000000000",
22107 => "0000000000000000",22108 => "0000000000000000",
22109 => "0000000000000000",22110 => "0000000000000000",
22111 => "0000000000000000",22112 => "0000000000000000",
22113 => "0000000000000000",22114 => "0000000000000000",
22115 => "0000000000000000",22116 => "0000000000000000",
22117 => "0000000000000000",22118 => "0000000000000000",
22119 => "0000000000000000",22120 => "0000000000000000",
22121 => "0000000000000000",22122 => "0000000000000000",
22123 => "0000000000000000",22124 => "0000000000000000",
22125 => "0000000000000000",22126 => "0000000000000000",
22127 => "0000000000000000",22128 => "0000000000000000",
22129 => "0000000000000000",22130 => "0000000000000000",
22131 => "0000000000000000",22132 => "0000000000000000",
22133 => "0000000000000000",22134 => "0000000000000000",
22135 => "0000000000000000",22136 => "0000000000000000",
22137 => "0000000000000000",22138 => "0000000000000000",
22139 => "0000000000000000",22140 => "0000000000000000",
22141 => "0000000000000000",22142 => "0000000000000000",
22143 => "0000000000000000",22144 => "0000000000000000",
22145 => "0000000000000000",22146 => "0000000000000000",
22147 => "0000000000000000",22148 => "0000000000000000",
22149 => "0000000000000000",22150 => "0000000000000000",
22151 => "0000000000000000",22152 => "0000000000000000",
22153 => "0000000000000000",22154 => "0000000000000000",
22155 => "0000000000000000",22156 => "0000000000000000",
22157 => "0000000000000000",22158 => "0000000000000000",
22159 => "0000000000000000",22160 => "0000000000000000",
22161 => "0000000000000000",22162 => "0000000000000000",
22163 => "0000000000000000",22164 => "0000000000000000",
22165 => "0000000000000000",22166 => "0000000000000000",
22167 => "0000000000000000",22168 => "0000000000000000",
22169 => "0000000000000000",22170 => "0000000000000000",
22171 => "0000000000000000",22172 => "0000000000000000",
22173 => "0000000000000000",22174 => "0000000000000000",
22175 => "0000000000000000",22176 => "0000000000000000",
22177 => "0000000000000000",22178 => "0000000000000000",
22179 => "0000000000000000",22180 => "0000000000000000",
22181 => "0000000000000000",22182 => "0000000000000000",
22183 => "0000000000000000",22184 => "0000000000000000",
22185 => "0000000000000000",22186 => "0000000000000000",
22187 => "0000000000000000",22188 => "0000000000000000",
22189 => "0000000000000000",22190 => "0000000000000000",
22191 => "0000000000000000",22192 => "0000000000000000",
22193 => "0000000000000000",22194 => "0000000000000000",
22195 => "0000000000000000",22196 => "0000000000000000",
22197 => "0000000000000000",22198 => "0000000000000000",
22199 => "0000000000000000",22200 => "0000000000000000",
22201 => "0000000000000000",22202 => "0000000000000000",
22203 => "0000000000000000",22204 => "0000000000000000",
22205 => "0000000000000000",22206 => "0000000000000000",
22207 => "0000000000000000",22208 => "0000000000000000",
22209 => "0000000000000000",22210 => "0000000000000000",
22211 => "0000000000000000",22212 => "0000000000000000",
22213 => "0000000000000000",22214 => "0000000000000000",
22215 => "0000000000000000",22216 => "0000000000000000",
22217 => "0000000000000000",22218 => "0000000000000000",
22219 => "0000000000000000",22220 => "0000000000000000",
22221 => "0000000000000000",22222 => "0000000000000000",
22223 => "0000000000000000",22224 => "0000000000000000",
22225 => "0000000000000000",22226 => "0000000000000000",
22227 => "0000000000000000",22228 => "0000000000000000",
22229 => "0000000000000000",22230 => "0000000000000000",
22231 => "0000000000000000",22232 => "0000000000000000",
22233 => "0000000000000000",22234 => "0000000000000000",
22235 => "0000000000000000",22236 => "0000000000000000",
22237 => "0000000000000000",22238 => "0000000000000000",
22239 => "0000000000000000",22240 => "0000000000000000",
22241 => "0000000000000000",22242 => "0000000000000000",
22243 => "0000000000000000",22244 => "0000000000000000",
22245 => "0000000000000000",22246 => "0000000000000000",
22247 => "0000000000000000",22248 => "0000000000000000",
22249 => "0000000000000000",22250 => "0000000000000000",
22251 => "0000000000000000",22252 => "0000000000000000",
22253 => "0000000000000000",22254 => "0000000000000000",
22255 => "0000000000000000",22256 => "0000000000000000",
22257 => "0000000000000000",22258 => "0000000000000000",
22259 => "0000000000000000",22260 => "0000000000000000",
22261 => "0000000000000000",22262 => "0000000000000000",
22263 => "0000000000000000",22264 => "0000000000000000",
22265 => "0000000000000000",22266 => "0000000000000000",
22267 => "0000000000000000",22268 => "0000000000000000",
22269 => "0000000000000000",22270 => "0000000000000000",
22271 => "0000000000000000",22272 => "0000000000000000",
22273 => "0000000000000000",22274 => "0000000000000000",
22275 => "0000000000000000",22276 => "0000000000000000",
22277 => "0000000000000000",22278 => "0000000000000000",
22279 => "0000000000000000",22280 => "0000000000000000",
22281 => "0000000000000000",22282 => "0000000000000000",
22283 => "0000000000000000",22284 => "0000000000000000",
22285 => "0000000000000000",22286 => "0000000000000000",
22287 => "0000000000000000",22288 => "0000000000000000",
22289 => "0000000000000000",22290 => "0000000000000000",
22291 => "0000000000000000",22292 => "0000000000000000",
22293 => "0000000000000000",22294 => "0000000000000000",
22295 => "0000000000000000",22296 => "0000000000000000",
22297 => "0000000000000000",22298 => "0000000000000000",
22299 => "0000000000000000",22300 => "0000000000000000",
22301 => "0000000000000000",22302 => "0000000000000000",
22303 => "0000000000000000",22304 => "0000000000000000",
22305 => "0000000000000000",22306 => "0000000000000000",
22307 => "0000000000000000",22308 => "0000000000000000",
22309 => "0000000000000000",22310 => "0000000000000000",
22311 => "0000000000000000",22312 => "0000000000000000",
22313 => "0000000000000000",22314 => "0000000000000000",
22315 => "0000000000000000",22316 => "0000000000000000",
22317 => "0000000000000000",22318 => "0000000000000000",
22319 => "0000000000000000",22320 => "0000000000000000",
22321 => "0000000000000000",22322 => "0000000000000000",
22323 => "0000000000000000",22324 => "0000000000000000",
22325 => "0000000000000000",22326 => "0000000000000000",
22327 => "0000000000000000",22328 => "0000000000000000",
22329 => "0000000000000000",22330 => "0000000000000000",
22331 => "0000000000000000",22332 => "0000000000000000",
22333 => "0000000000000000",22334 => "0000000000000000",
22335 => "0000000000000000",22336 => "0000000000000000",
22337 => "0000000000000000",22338 => "0000000000000000",
22339 => "0000000000000000",22340 => "0000000000000000",
22341 => "0000000000000000",22342 => "0000000000000000",
22343 => "0000000000000000",22344 => "0000000000000000",
22345 => "0000000000000000",22346 => "0000000000000000",
22347 => "0000000000000000",22348 => "0000000000000000",
22349 => "0000000000000000",22350 => "0000000000000000",
22351 => "0000000000000000",22352 => "0000000000000000",
22353 => "0000000000000000",22354 => "0000000000000000",
22355 => "0000000000000000",22356 => "0000000000000000",
22357 => "0000000000000000",22358 => "0000000000000000",
22359 => "0000000000000000",22360 => "0000000000000000",
22361 => "0000000000000000",22362 => "0000000000000000",
22363 => "0000000000000000",22364 => "0000000000000000",
22365 => "0000000000000000",22366 => "0000000000000000",
22367 => "0000000000000000",22368 => "0000000000000000",
22369 => "0000000000000000",22370 => "0000000000000000",
22371 => "0000000000000000",22372 => "0000000000000000",
22373 => "0000000000000000",22374 => "0000000000000000",
22375 => "0000000000000000",22376 => "0000000000000000",
22377 => "0000000000000000",22378 => "0000000000000000",
22379 => "0000000000000000",22380 => "0000000000000000",
22381 => "0000000000000000",22382 => "0000000000000000",
22383 => "0000000000000000",22384 => "0000000000000000",
22385 => "0000000000000000",22386 => "0000000000000000",
22387 => "0000000000000000",22388 => "0000000000000000",
22389 => "0000000000000000",22390 => "0000000000000000",
22391 => "0000000000000000",22392 => "0000000000000000",
22393 => "0000000000000000",22394 => "0000000000000000",
22395 => "0000000000000000",22396 => "0000000000000000",
22397 => "0000000000000000",22398 => "0000000000000000",
22399 => "0000000000000000",22400 => "0000000000000000",
22401 => "0000000000000000",22402 => "0000000000000000",
22403 => "0000000000000000",22404 => "0000000000000000",
22405 => "0000000000000000",22406 => "0000000000000000",
22407 => "0000000000000000",22408 => "0000000000000000",
22409 => "0000000000000000",22410 => "0000000000000000",
22411 => "0000000000000000",22412 => "0000000000000000",
22413 => "0000000000000000",22414 => "0000000000000000",
22415 => "0000000000000000",22416 => "0000000000000000",
22417 => "0000000000000000",22418 => "0000000000000000",
22419 => "0000000000000000",22420 => "0000000000000000",
22421 => "0000000000000000",22422 => "0000000000000000",
22423 => "0000000000000000",22424 => "0000000000000000",
22425 => "0000000000000000",22426 => "0000000000000000",
22427 => "0000000000000000",22428 => "0000000000000000",
22429 => "0000000000000000",22430 => "0000000000000000",
22431 => "0000000000000000",22432 => "0000000000000000",
22433 => "0000000000000000",22434 => "0000000000000000",
22435 => "0000000000000000",22436 => "0000000000000000",
22437 => "0000000000000000",22438 => "0000000000000000",
22439 => "0000000000000000",22440 => "0000000000000000",
22441 => "0000000000000000",22442 => "0000000000000000",
22443 => "0000000000000000",22444 => "0000000000000000",
22445 => "0000000000000000",22446 => "0000000000000000",
22447 => "0000000000000000",22448 => "0000000000000000",
22449 => "0000000000000000",22450 => "0000000000000000",
22451 => "0000000000000000",22452 => "0000000000000000",
22453 => "0000000000000000",22454 => "0000000000000000",
22455 => "0000000000000000",22456 => "0000000000000000",
22457 => "0000000000000000",22458 => "0000000000000000",
22459 => "0000000000000000",22460 => "0000000000000000",
22461 => "0000000000000000",22462 => "0000000000000000",
22463 => "0000000000000000",22464 => "0000000000000000",
22465 => "0000000000000000",22466 => "0000000000000000",
22467 => "0000000000000000",22468 => "0000000000000000",
22469 => "0000000000000000",22470 => "0000000000000000",
22471 => "0000000000000000",22472 => "0000000000000000",
22473 => "0000000000000000",22474 => "0000000000000000",
22475 => "0000000000000000",22476 => "0000000000000000",
22477 => "0000000000000000",22478 => "0000000000000000",
22479 => "0000000000000000",22480 => "0000000000000000",
22481 => "0000000000000000",22482 => "0000000000000000",
22483 => "0000000000000000",22484 => "0000000000000000",
22485 => "0000000000000000",22486 => "0000000000000000",
22487 => "0000000000000000",22488 => "0000000000000000",
22489 => "0000000000000000",22490 => "0000000000000000",
22491 => "0000000000000000",22492 => "0000000000000000",
22493 => "0000000000000000",22494 => "0000000000000000",
22495 => "0000000000000000",22496 => "0000000000000000",
22497 => "0000000000000000",22498 => "0000000000000000",
22499 => "0000000000000000",22500 => "0000000000000000",
22501 => "0000000000000000",22502 => "0000000000000000",
22503 => "0000000000000000",22504 => "0000000000000000",
22505 => "0000000000000000",22506 => "0000000000000000",
22507 => "0000000000000000",22508 => "0000000000000000",
22509 => "0000000000000000",22510 => "0000000000000000",
22511 => "0000000000000000",22512 => "0000000000000000",
22513 => "0000000000000000",22514 => "0000000000000000",
22515 => "0000000000000000",22516 => "0000000000000000",
22517 => "0000000000000000",22518 => "0000000000000000",
22519 => "0000000000000000",22520 => "0000000000000000",
22521 => "0000000000000000",22522 => "0000000000000000",
22523 => "0000000000000000",22524 => "0000000000000000",
22525 => "0000000000000000",22526 => "0000000000000000",
22527 => "0000000000000000",22528 => "0000000000000000",
22529 => "0000000000000000",22530 => "0000000000000000",
22531 => "0000000000000000",22532 => "0000000000000000",
22533 => "0000000000000000",22534 => "0000000000000000",
22535 => "0000000000000000",22536 => "0000000000000000",
22537 => "0000000000000000",22538 => "0000000000000000",
22539 => "0000000000000000",22540 => "0000000000000000",
22541 => "0000000000000000",22542 => "0000000000000000",
22543 => "0000000000000000",22544 => "0000000000000000",
22545 => "0000000000000000",22546 => "0000000000000000",
22547 => "0000000000000000",22548 => "0000000000000000",
22549 => "0000000000000000",22550 => "0000000000000000",
22551 => "0000000000000000",22552 => "0000000000000000",
22553 => "0000000000000000",22554 => "0000000000000000",
22555 => "0000000000000000",22556 => "0000000000000000",
22557 => "0000000000000000",22558 => "0000000000000000",
22559 => "0000000000000000",22560 => "0000000000000000",
22561 => "0000000000000000",22562 => "0000000000000000",
22563 => "0000000000000000",22564 => "0000000000000000",
22565 => "0000000000000000",22566 => "0000000000000000",
22567 => "0000000000000000",22568 => "0000000000000000",
22569 => "0000000000000000",22570 => "0000000000000000",
22571 => "0000000000000000",22572 => "0000000000000000",
22573 => "0000000000000000",22574 => "0000000000000000",
22575 => "0000000000000000",22576 => "0000000000000000",
22577 => "0000000000000000",22578 => "0000000000000000",
22579 => "0000000000000000",22580 => "0000000000000000",
22581 => "0000000000000000",22582 => "0000000000000000",
22583 => "0000000000000000",22584 => "0000000000000000",
22585 => "0000000000000000",22586 => "0000000000000000",
22587 => "0000000000000000",22588 => "0000000000000000",
22589 => "0000000000000000",22590 => "0000000000000000",
22591 => "0000000000000000",22592 => "0000000000000000",
22593 => "0000000000000000",22594 => "0000000000000000",
22595 => "0000000000000000",22596 => "0000000000000000",
22597 => "0000000000000000",22598 => "0000000000000000",
22599 => "0000000000000000",22600 => "0000000000000000",
22601 => "0000000000000000",22602 => "0000000000000000",
22603 => "0000000000000000",22604 => "0000000000000000",
22605 => "0000000000000000",22606 => "0000000000000000",
22607 => "0000000000000000",22608 => "0000000000000000",
22609 => "0000000000000000",22610 => "0000000000000000",
22611 => "0000000000000000",22612 => "0000000000000000",
22613 => "0000000000000000",22614 => "0000000000000000",
22615 => "0000000000000000",22616 => "0000000000000000",
22617 => "0000000000000000",22618 => "0000000000000000",
22619 => "0000000000000000",22620 => "0000000000000000",
22621 => "0000000000000000",22622 => "0000000000000000",
22623 => "0000000000000000",22624 => "0000000000000000",
22625 => "0000000000000000",22626 => "0000000000000000",
22627 => "0000000000000000",22628 => "0000000000000000",
22629 => "0000000000000000",22630 => "0000000000000000",
22631 => "0000000000000000",22632 => "0000000000000000",
22633 => "0000000000000000",22634 => "0000000000000000",
22635 => "0000000000000000",22636 => "0000000000000000",
22637 => "0000000000000000",22638 => "0000000000000000",
22639 => "0000000000000000",22640 => "0000000000000000",
22641 => "0000000000000000",22642 => "0000000000000000",
22643 => "0000000000000000",22644 => "0000000000000000",
22645 => "0000000000000000",22646 => "0000000000000000",
22647 => "0000000000000000",22648 => "0000000000000000",
22649 => "0000000000000000",22650 => "0000000000000000",
22651 => "0000000000000000",22652 => "0000000000000000",
22653 => "0000000000000000",22654 => "0000000000000000",
22655 => "0000000000000000",22656 => "0000000000000000",
22657 => "0000000000000000",22658 => "0000000000000000",
22659 => "0000000000000000",22660 => "0000000000000000",
22661 => "0000000000000000",22662 => "0000000000000000",
22663 => "0000000000000000",22664 => "0000000000000000",
22665 => "0000000000000000",22666 => "0000000000000000",
22667 => "0000000000000000",22668 => "0000000000000000",
22669 => "0000000000000000",22670 => "0000000000000000",
22671 => "0000000000000000",22672 => "0000000000000000",
22673 => "0000000000000000",22674 => "0000000000000000",
22675 => "0000000000000000",22676 => "0000000000000000",
22677 => "0000000000000000",22678 => "0000000000000000",
22679 => "0000000000000000",22680 => "0000000000000000",
22681 => "0000000000000000",22682 => "0000000000000000",
22683 => "0000000000000000",22684 => "0000000000000000",
22685 => "0000000000000000",22686 => "0000000000000000",
22687 => "0000000000000000",22688 => "0000000000000000",
22689 => "0000000000000000",22690 => "0000000000000000",
22691 => "0000000000000000",22692 => "0000000000000000",
22693 => "0000000000000000",22694 => "0000000000000000",
22695 => "0000000000000000",22696 => "0000000000000000",
22697 => "0000000000000000",22698 => "0000000000000000",
22699 => "0000000000000000",22700 => "0000000000000000",
22701 => "0000000000000000",22702 => "0000000000000000",
22703 => "0000000000000000",22704 => "0000000000000000",
22705 => "0000000000000000",22706 => "0000000000000000",
22707 => "0000000000000000",22708 => "0000000000000000",
22709 => "0000000000000000",22710 => "0000000000000000",
22711 => "0000000000000000",22712 => "0000000000000000",
22713 => "0000000000000000",22714 => "0000000000000000",
22715 => "0000000000000000",22716 => "0000000000000000",
22717 => "0000000000000000",22718 => "0000000000000000",
22719 => "0000000000000000",22720 => "0000000000000000",
22721 => "0000000000000000",22722 => "0000000000000000",
22723 => "0000000000000000",22724 => "0000000000000000",
22725 => "0000000000000000",22726 => "0000000000000000",
22727 => "0000000000000000",22728 => "0000000000000000",
22729 => "0000000000000000",22730 => "0000000000000000",
22731 => "0000000000000000",22732 => "0000000000000000",
22733 => "0000000000000000",22734 => "0000000000000000",
22735 => "0000000000000000",22736 => "0000000000000000",
22737 => "0000000000000000",22738 => "0000000000000000",
22739 => "0000000000000000",22740 => "0000000000000000",
22741 => "0000000000000000",22742 => "0000000000000000",
22743 => "0000000000000000",22744 => "0000000000000000",
22745 => "0000000000000000",22746 => "0000000000000000",
22747 => "0000000000000000",22748 => "0000000000000000",
22749 => "0000000000000000",22750 => "0000000000000000",
22751 => "0000000000000000",22752 => "0000000000000000",
22753 => "0000000000000000",22754 => "0000000000000000",
22755 => "0000000000000000",22756 => "0000000000000000",
22757 => "0000000000000000",22758 => "0000000000000000",
22759 => "0000000000000000",22760 => "0000000000000000",
22761 => "0000000000000000",22762 => "0000000000000000",
22763 => "0000000000000000",22764 => "0000000000000000",
22765 => "0000000000000000",22766 => "0000000000000000",
22767 => "0000000000000000",22768 => "0000000000000000",
22769 => "0000000000000000",22770 => "0000000000000000",
22771 => "0000000000000000",22772 => "0000000000000000",
22773 => "0000000000000000",22774 => "0000000000000000",
22775 => "0000000000000000",22776 => "0000000000000000",
22777 => "0000000000000000",22778 => "0000000000000000",
22779 => "0000000000000000",22780 => "0000000000000000",
22781 => "0000000000000000",22782 => "0000000000000000",
22783 => "0000000000000000",22784 => "0000000000000000",
22785 => "0000000000000000",22786 => "0000000000000000",
22787 => "0000000000000000",22788 => "0000000000000000",
22789 => "0000000000000000",22790 => "0000000000000000",
22791 => "0000000000000000",22792 => "0000000000000000",
22793 => "0000000000000000",22794 => "0000000000000000",
22795 => "0000000000000000",22796 => "0000000000000000",
22797 => "0000000000000000",22798 => "0000000000000000",
22799 => "0000000000000000",22800 => "0000000000000000",
22801 => "0000000000000000",22802 => "0000000000000000",
22803 => "0000000000000000",22804 => "0000000000000000",
22805 => "0000000000000000",22806 => "0000000000000000",
22807 => "0000000000000000",22808 => "0000000000000000",
22809 => "0000000000000000",22810 => "0000000000000000",
22811 => "0000000000000000",22812 => "0000000000000000",
22813 => "0000000000000000",22814 => "0000000000000000",
22815 => "0000000000000000",22816 => "0000000000000000",
22817 => "0000000000000000",22818 => "0000000000000000",
22819 => "0000000000000000",22820 => "0000000000000000",
22821 => "0000000000000000",22822 => "0000000000000000",
22823 => "0000000000000000",22824 => "0000000000000000",
22825 => "0000000000000000",22826 => "0000000000000000",
22827 => "0000000000000000",22828 => "0000000000000000",
22829 => "0000000000000000",22830 => "0000000000000000",
22831 => "0000000000000000",22832 => "0000000000000000",
22833 => "0000000000000000",22834 => "0000000000000000",
22835 => "0000000000000000",22836 => "0000000000000000",
22837 => "0000000000000000",22838 => "0000000000000000",
22839 => "0000000000000000",22840 => "0000000000000000",
22841 => "0000000000000000",22842 => "0000000000000000",
22843 => "0000000000000000",22844 => "0000000000000000",
22845 => "0000000000000000",22846 => "0000000000000000",
22847 => "0000000000000000",22848 => "0000000000000000",
22849 => "0000000000000000",22850 => "0000000000000000",
22851 => "0000000000000000",22852 => "0000000000000000",
22853 => "0000000000000000",22854 => "0000000000000000",
22855 => "0000000000000000",22856 => "0000000000000000",
22857 => "0000000000000000",22858 => "0000000000000000",
22859 => "0000000000000000",22860 => "0000000000000000",
22861 => "0000000000000000",22862 => "0000000000000000",
22863 => "0000000000000000",22864 => "0000000000000000",
22865 => "0000000000000000",22866 => "0000000000000000",
22867 => "0000000000000000",22868 => "0000000000000000",
22869 => "0000000000000000",22870 => "0000000000000000",
22871 => "0000000000000000",22872 => "0000000000000000",
22873 => "0000000000000000",22874 => "0000000000000000",
22875 => "0000000000000000",22876 => "0000000000000000",
22877 => "0000000000000000",22878 => "0000000000000000",
22879 => "0000000000000000",22880 => "0000000000000000",
22881 => "0000000000000000",22882 => "0000000000000000",
22883 => "0000000000000000",22884 => "0000000000000000",
22885 => "0000000000000000",22886 => "0000000000000000",
22887 => "0000000000000000",22888 => "0000000000000000",
22889 => "0000000000000000",22890 => "0000000000000000",
22891 => "0000000000000000",22892 => "0000000000000000",
22893 => "0000000000000000",22894 => "0000000000000000",
22895 => "0000000000000000",22896 => "0000000000000000",
22897 => "0000000000000000",22898 => "0000000000000000",
22899 => "0000000000000000",22900 => "0000000000000000",
22901 => "0000000000000000",22902 => "0000000000000000",
22903 => "0000000000000000",22904 => "0000000000000000",
22905 => "0000000000000000",22906 => "0000000000000000",
22907 => "0000000000000000",22908 => "0000000000000000",
22909 => "0000000000000000",22910 => "0000000000000000",
22911 => "0000000000000000",22912 => "0000000000000000",
22913 => "0000000000000000",22914 => "0000000000000000",
22915 => "0000000000000000",22916 => "0000000000000000",
22917 => "0000000000000000",22918 => "0000000000000000",
22919 => "0000000000000000",22920 => "0000000000000000",
22921 => "0000000000000000",22922 => "0000000000000000",
22923 => "0000000000000000",22924 => "0000000000000000",
22925 => "0000000000000000",22926 => "0000000000000000",
22927 => "0000000000000000",22928 => "0000000000000000",
22929 => "0000000000000000",22930 => "0000000000000000",
22931 => "0000000000000000",22932 => "0000000000000000",
22933 => "0000000000000000",22934 => "0000000000000000",
22935 => "0000000000000000",22936 => "0000000000000000",
22937 => "0000000000000000",22938 => "0000000000000000",
22939 => "0000000000000000",22940 => "0000000000000000",
22941 => "0000000000000000",22942 => "0000000000000000",
22943 => "0000000000000000",22944 => "0000000000000000",
22945 => "0000000000000000",22946 => "0000000000000000",
22947 => "0000000000000000",22948 => "0000000000000000",
22949 => "0000000000000000",22950 => "0000000000000000",
22951 => "0000000000000000",22952 => "0000000000000000",
22953 => "0000000000000000",22954 => "0000000000000000",
22955 => "0000000000000000",22956 => "0000000000000000",
22957 => "0000000000000000",22958 => "0000000000000000",
22959 => "0000000000000000",22960 => "0000000000000000",
22961 => "0000000000000000",22962 => "0000000000000000",
22963 => "0000000000000000",22964 => "0000000000000000",
22965 => "0000000000000000",22966 => "0000000000000000",
22967 => "0000000000000000",22968 => "0000000000000000",
22969 => "0000000000000000",22970 => "0000000000000000",
22971 => "0000000000000000",22972 => "0000000000000000",
22973 => "0000000000000000",22974 => "0000000000000000",
22975 => "0000000000000000",22976 => "0000000000000000",
22977 => "0000000000000000",22978 => "0000000000000000",
22979 => "0000000000000000",22980 => "0000000000000000",
22981 => "0000000000000000",22982 => "0000000000000000",
22983 => "0000000000000000",22984 => "0000000000000000",
22985 => "0000000000000000",22986 => "0000000000000000",
22987 => "0000000000000000",22988 => "0000000000000000",
22989 => "0000000000000000",22990 => "0000000000000000",
22991 => "0000000000000000",22992 => "0000000000000000",
22993 => "0000000000000000",22994 => "0000000000000000",
22995 => "0000000000000000",22996 => "0000000000000000",
22997 => "0000000000000000",22998 => "0000000000000000",
22999 => "0000000000000000",23000 => "0000000000000000",
23001 => "0000000000000000",23002 => "0000000000000000",
23003 => "0000000000000000",23004 => "0000000000000000",
23005 => "0000000000000000",23006 => "0000000000000000",
23007 => "0000000000000000",23008 => "0000000000000000",
23009 => "0000000000000000",23010 => "0000000000000000",
23011 => "0000000000000000",23012 => "0000000000000000",
23013 => "0000000000000000",23014 => "0000000000000000",
23015 => "0000000000000000",23016 => "0000000000000000",
23017 => "0000000000000000",23018 => "0000000000000000",
23019 => "0000000000000000",23020 => "0000000000000000",
23021 => "0000000000000000",23022 => "0000000000000000",
23023 => "0000000000000000",23024 => "0000000000000000",
23025 => "0000000000000000",23026 => "0000000000000000",
23027 => "0000000000000000",23028 => "0000000000000000",
23029 => "0000000000000000",23030 => "0000000000000000",
23031 => "0000000000000000",23032 => "0000000000000000",
23033 => "0000000000000000",23034 => "0000000000000000",
23035 => "0000000000000000",23036 => "0000000000000000",
23037 => "0000000000000000",23038 => "0000000000000000",
23039 => "0000000000000000",23040 => "0000000000000000",
23041 => "0000000000000000",23042 => "0000000000000000",
23043 => "0000000000000000",23044 => "0000000000000000",
23045 => "0000000000000000",23046 => "0000000000000000",
23047 => "0000000000000000",23048 => "0000000000000000",
23049 => "0000000000000000",23050 => "0000000000000000",
23051 => "0000000000000000",23052 => "0000000000000000",
23053 => "0000000000000000",23054 => "0000000000000000",
23055 => "0000000000000000",23056 => "0000000000000000",
23057 => "0000000000000000",23058 => "0000000000000000",
23059 => "0000000000000000",23060 => "0000000000000000",
23061 => "0000000000000000",23062 => "0000000000000000",
23063 => "0000000000000000",23064 => "0000000000000000",
23065 => "0000000000000000",23066 => "0000000000000000",
23067 => "0000000000000000",23068 => "0000000000000000",
23069 => "0000000000000000",23070 => "0000000000000000",
23071 => "0000000000000000",23072 => "0000000000000000",
23073 => "0000000000000000",23074 => "0000000000000000",
23075 => "0000000000000000",23076 => "0000000000000000",
23077 => "0000000000000000",23078 => "0000000000000000",
23079 => "0000000000000000",23080 => "0000000000000000",
23081 => "0000000000000000",23082 => "0000000000000000",
23083 => "0000000000000000",23084 => "0000000000000000",
23085 => "0000000000000000",23086 => "0000000000000000",
23087 => "0000000000000000",23088 => "0000000000000000",
23089 => "0000000000000000",23090 => "0000000000000000",
23091 => "0000000000000000",23092 => "0000000000000000",
23093 => "0000000000000000",23094 => "0000000000000000",
23095 => "0000000000000000",23096 => "0000000000000000",
23097 => "0000000000000000",23098 => "0000000000000000",
23099 => "0000000000000000",23100 => "0000000000000000",
23101 => "0000000000000000",23102 => "0000000000000000",
23103 => "0000000000000000",23104 => "0000000000000000",
23105 => "0000000000000000",23106 => "0000000000000000",
23107 => "0000000000000000",23108 => "0000000000000000",
23109 => "0000000000000000",23110 => "0000000000000000",
23111 => "0000000000000000",23112 => "0000000000000000",
23113 => "0000000000000000",23114 => "0000000000000000",
23115 => "0000000000000000",23116 => "0000000000000000",
23117 => "0000000000000000",23118 => "0000000000000000",
23119 => "0000000000000000",23120 => "0000000000000000",
23121 => "0000000000000000",23122 => "0000000000000000",
23123 => "0000000000000000",23124 => "0000000000000000",
23125 => "0000000000000000",23126 => "0000000000000000",
23127 => "0000000000000000",23128 => "0000000000000000",
23129 => "0000000000000000",23130 => "0000000000000000",
23131 => "0000000000000000",23132 => "0000000000000000",
23133 => "0000000000000000",23134 => "0000000000000000",
23135 => "0000000000000000",23136 => "0000000000000000",
23137 => "0000000000000000",23138 => "0000000000000000",
23139 => "0000000000000000",23140 => "0000000000000000",
23141 => "0000000000000000",23142 => "0000000000000000",
23143 => "0000000000000000",23144 => "0000000000000000",
23145 => "0000000000000000",23146 => "0000000000000000",
23147 => "0000000000000000",23148 => "0000000000000000",
23149 => "0000000000000000",23150 => "0000000000000000",
23151 => "0000000000000000",23152 => "0000000000000000",
23153 => "0000000000000000",23154 => "0000000000000000",
23155 => "0000000000000000",23156 => "0000000000000000",
23157 => "0000000000000000",23158 => "0000000000000000",
23159 => "0000000000000000",23160 => "0000000000000000",
23161 => "0000000000000000",23162 => "0000000000000000",
23163 => "0000000000000000",23164 => "0000000000000000",
23165 => "0000000000000000",23166 => "0000000000000000",
23167 => "0000000000000000",23168 => "0000000000000000",
23169 => "0000000000000000",23170 => "0000000000000000",
23171 => "0000000000000000",23172 => "0000000000000000",
23173 => "0000000000000000",23174 => "0000000000000000",
23175 => "0000000000000000",23176 => "0000000000000000",
23177 => "0000000000000000",23178 => "0000000000000000",
23179 => "0000000000000000",23180 => "0000000000000000",
23181 => "0000000000000000",23182 => "0000000000000000",
23183 => "0000000000000000",23184 => "0000000000000000",
23185 => "0000000000000000",23186 => "0000000000000000",
23187 => "0000000000000000",23188 => "0000000000000000",
23189 => "0000000000000000",23190 => "0000000000000000",
23191 => "0000000000000000",23192 => "0000000000000000",
23193 => "0000000000000000",23194 => "0000000000000000",
23195 => "0000000000000000",23196 => "0000000000000000",
23197 => "0000000000000000",23198 => "0000000000000000",
23199 => "0000000000000000",23200 => "0000000000000000",
23201 => "0000000000000000",23202 => "0000000000000000",
23203 => "0000000000000000",23204 => "0000000000000000",
23205 => "0000000000000000",23206 => "0000000000000000",
23207 => "0000000000000000",23208 => "0000000000000000",
23209 => "0000000000000000",23210 => "0000000000000000",
23211 => "0000000000000000",23212 => "0000000000000000",
23213 => "0000000000000000",23214 => "0000000000000000",
23215 => "0000000000000000",23216 => "0000000000000000",
23217 => "0000000000000000",23218 => "0000000000000000",
23219 => "0000000000000000",23220 => "0000000000000000",
23221 => "0000000000000000",23222 => "0000000000000000",
23223 => "0000000000000000",23224 => "0000000000000000",
23225 => "0000000000000000",23226 => "0000000000000000",
23227 => "0000000000000000",23228 => "0000000000000000",
23229 => "0000000000000000",23230 => "0000000000000000",
23231 => "0000000000000000",23232 => "0000000000000000",
23233 => "0000000000000000",23234 => "0000000000000000",
23235 => "0000000000000000",23236 => "0000000000000000",
23237 => "0000000000000000",23238 => "0000000000000000",
23239 => "0000000000000000",23240 => "0000000000000000",
23241 => "0000000000000000",23242 => "0000000000000000",
23243 => "0000000000000000",23244 => "0000000000000000",
23245 => "0000000000000000",23246 => "0000000000000000",
23247 => "0000000000000000",23248 => "0000000000000000",
23249 => "0000000000000000",23250 => "0000000000000000",
23251 => "0000000000000000",23252 => "0000000000000000",
23253 => "0000000000000000",23254 => "0000000000000000",
23255 => "0000000000000000",23256 => "0000000000000000",
23257 => "0000000000000000",23258 => "0000000000000000",
23259 => "0000000000000000",23260 => "0000000000000000",
23261 => "0000000000000000",23262 => "0000000000000000",
23263 => "0000000000000000",23264 => "0000000000000000",
23265 => "0000000000000000",23266 => "0000000000000000",
23267 => "0000000000000000",23268 => "0000000000000000",
23269 => "0000000000000000",23270 => "0000000000000000",
23271 => "0000000000000000",23272 => "0000000000000000",
23273 => "0000000000000000",23274 => "0000000000000000",
23275 => "0000000000000000",23276 => "0000000000000000",
23277 => "0000000000000000",23278 => "0000000000000000",
23279 => "0000000000000000",23280 => "0000000000000000",
23281 => "0000000000000000",23282 => "0000000000000000",
23283 => "0000000000000000",23284 => "0000000000000000",
23285 => "0000000000000000",23286 => "0000000000000000",
23287 => "0000000000000000",23288 => "0000000000000000",
23289 => "0000000000000000",23290 => "0000000000000000",
23291 => "0000000000000000",23292 => "0000000000000000",
23293 => "0000000000000000",23294 => "0000000000000000",
23295 => "0000000000000000",23296 => "0000000000000000",
23297 => "0000000000000000",23298 => "0000000000000000",
23299 => "0000000000000000",23300 => "0000000000000000",
23301 => "0000000000000000",23302 => "0000000000000000",
23303 => "0000000000000000",23304 => "0000000000000000",
23305 => "0000000000000000",23306 => "0000000000000000",
23307 => "0000000000000000",23308 => "0000000000000000",
23309 => "0000000000000000",23310 => "0000000000000000",
23311 => "0000000000000000",23312 => "0000000000000000",
23313 => "0000000000000000",23314 => "0000000000000000",
23315 => "0000000000000000",23316 => "0000000000000000",
23317 => "0000000000000000",23318 => "0000000000000000",
23319 => "0000000000000000",23320 => "0000000000000000",
23321 => "0000000000000000",23322 => "0000000000000000",
23323 => "0000000000000000",23324 => "0000000000000000",
23325 => "0000000000000000",23326 => "0000000000000000",
23327 => "0000000000000000",23328 => "0000000000000000",
23329 => "0000000000000000",23330 => "0000000000000000",
23331 => "0000000000000000",23332 => "0000000000000000",
23333 => "0000000000000000",23334 => "0000000000000000",
23335 => "0000000000000000",23336 => "0000000000000000",
23337 => "0000000000000000",23338 => "0000000000000000",
23339 => "0000000000000000",23340 => "0000000000000000",
23341 => "0000000000000000",23342 => "0000000000000000",
23343 => "0000000000000000",23344 => "0000000000000000",
23345 => "0000000000000000",23346 => "0000000000000000",
23347 => "0000000000000000",23348 => "0000000000000000",
23349 => "0000000000000000",23350 => "0000000000000000",
23351 => "0000000000000000",23352 => "0000000000000000",
23353 => "0000000000000000",23354 => "0000000000000000",
23355 => "0000000000000000",23356 => "0000000000000000",
23357 => "0000000000000000",23358 => "0000000000000000",
23359 => "0000000000000000",23360 => "0000000000000000",
23361 => "0000000000000000",23362 => "0000000000000000",
23363 => "0000000000000000",23364 => "0000000000000000",
23365 => "0000000000000000",23366 => "0000000000000000",
23367 => "0000000000000000",23368 => "0000000000000000",
23369 => "0000000000000000",23370 => "0000000000000000",
23371 => "0000000000000000",23372 => "0000000000000000",
23373 => "0000000000000000",23374 => "0000000000000000",
23375 => "0000000000000000",23376 => "0000000000000000",
23377 => "0000000000000000",23378 => "0000000000000000",
23379 => "0000000000000000",23380 => "0000000000000000",
23381 => "0000000000000000",23382 => "0000000000000000",
23383 => "0000000000000000",23384 => "0000000000000000",
23385 => "0000000000000000",23386 => "0000000000000000",
23387 => "0000000000000000",23388 => "0000000000000000",
23389 => "0000000000000000",23390 => "0000000000000000",
23391 => "0000000000000000",23392 => "0000000000000000",
23393 => "0000000000000000",23394 => "0000000000000000",
23395 => "0000000000000000",23396 => "0000000000000000",
23397 => "0000000000000000",23398 => "0000000000000000",
23399 => "0000000000000000",23400 => "0000000000000000",
23401 => "0000000000000000",23402 => "0000000000000000",
23403 => "0000000000000000",23404 => "0000000000000000",
23405 => "0000000000000000",23406 => "0000000000000000",
23407 => "0000000000000000",23408 => "0000000000000000",
23409 => "0000000000000000",23410 => "0000000000000000",
23411 => "0000000000000000",23412 => "0000000000000000",
23413 => "0000000000000000",23414 => "0000000000000000",
23415 => "0000000000000000",23416 => "0000000000000000",
23417 => "0000000000000000",23418 => "0000000000000000",
23419 => "0000000000000000",23420 => "0000000000000000",
23421 => "0000000000000000",23422 => "0000000000000000",
23423 => "0000000000000000",23424 => "0000000000000000",
23425 => "0000000000000000",23426 => "0000000000000000",
23427 => "0000000000000000",23428 => "0000000000000000",
23429 => "0000000000000000",23430 => "0000000000000000",
23431 => "0000000000000000",23432 => "0000000000000000",
23433 => "0000000000000000",23434 => "0000000000000000",
23435 => "0000000000000000",23436 => "0000000000000000",
23437 => "0000000000000000",23438 => "0000000000000000",
23439 => "0000000000000000",23440 => "0000000000000000",
23441 => "0000000000000000",23442 => "0000000000000000",
23443 => "0000000000000000",23444 => "0000000000000000",
23445 => "0000000000000000",23446 => "0000000000000000",
23447 => "0000000000000000",23448 => "0000000000000000",
23449 => "0000000000000000",23450 => "0000000000000000",
23451 => "0000000000000000",23452 => "0000000000000000",
23453 => "0000000000000000",23454 => "0000000000000000",
23455 => "0000000000000000",23456 => "0000000000000000",
23457 => "0000000000000000",23458 => "0000000000000000",
23459 => "0000000000000000",23460 => "0000000000000000",
23461 => "0000000000000000",23462 => "0000000000000000",
23463 => "0000000000000000",23464 => "0000000000000000",
23465 => "0000000000000000",23466 => "0000000000000000",
23467 => "0000000000000000",23468 => "0000000000000000",
23469 => "0000000000000000",23470 => "0000000000000000",
23471 => "0000000000000000",23472 => "0000000000000000",
23473 => "0000000000000000",23474 => "0000000000000000",
23475 => "0000000000000000",23476 => "0000000000000000",
23477 => "0000000000000000",23478 => "0000000000000000",
23479 => "0000000000000000",23480 => "0000000000000000",
23481 => "0000000000000000",23482 => "0000000000000000",
23483 => "0000000000000000",23484 => "0000000000000000",
23485 => "0000000000000000",23486 => "0000000000000000",
23487 => "0000000000000000",23488 => "0000000000000000",
23489 => "0000000000000000",23490 => "0000000000000000",
23491 => "0000000000000000",23492 => "0000000000000000",
23493 => "0000000000000000",23494 => "0000000000000000",
23495 => "0000000000000000",23496 => "0000000000000000",
23497 => "0000000000000000",23498 => "0000000000000000",
23499 => "0000000000000000",23500 => "0000000000000000",
23501 => "0000000000000000",23502 => "0000000000000000",
23503 => "0000000000000000",23504 => "0000000000000000",
23505 => "0000000000000000",23506 => "0000000000000000",
23507 => "0000000000000000",23508 => "0000000000000000",
23509 => "0000000000000000",23510 => "0000000000000000",
23511 => "0000000000000000",23512 => "0000000000000000",
23513 => "0000000000000000",23514 => "0000000000000000",
23515 => "0000000000000000",23516 => "0000000000000000",
23517 => "0000000000000000",23518 => "0000000000000000",
23519 => "0000000000000000",23520 => "0000000000000000",
23521 => "0000000000000000",23522 => "0000000000000000",
23523 => "0000000000000000",23524 => "0000000000000000",
23525 => "0000000000000000",23526 => "0000000000000000",
23527 => "0000000000000000",23528 => "0000000000000000",
23529 => "0000000000000000",23530 => "0000000000000000",
23531 => "0000000000000000",23532 => "0000000000000000",
23533 => "0000000000000000",23534 => "0000000000000000",
23535 => "0000000000000000",23536 => "0000000000000000",
23537 => "0000000000000000",23538 => "0000000000000000",
23539 => "0000000000000000",23540 => "0000000000000000",
23541 => "0000000000000000",23542 => "0000000000000000",
23543 => "0000000000000000",23544 => "0000000000000000",
23545 => "0000000000000000",23546 => "0000000000000000",
23547 => "0000000000000000",23548 => "0000000000000000",
23549 => "0000000000000000",23550 => "0000000000000000",
23551 => "0000000000000000",23552 => "0000000000000000",
23553 => "0000000000000000",23554 => "0000000000000000",
23555 => "0000000000000000",23556 => "0000000000000000",
23557 => "0000000000000000",23558 => "0000000000000000",
23559 => "0000000000000000",23560 => "0000000000000000",
23561 => "0000000000000000",23562 => "0000000000000000",
23563 => "0000000000000000",23564 => "0000000000000000",
23565 => "0000000000000000",23566 => "0000000000000000",
23567 => "0000000000000000",23568 => "0000000000000000",
23569 => "0000000000000000",23570 => "0000000000000000",
23571 => "0000000000000000",23572 => "0000000000000000",
23573 => "0000000000000000",23574 => "0000000000000000",
23575 => "0000000000000000",23576 => "0000000000000000",
23577 => "0000000000000000",23578 => "0000000000000000",
23579 => "0000000000000000",23580 => "0000000000000000",
23581 => "0000000000000000",23582 => "0000000000000000",
23583 => "0000000000000000",23584 => "0000000000000000",
23585 => "0000000000000000",23586 => "0000000000000000",
23587 => "0000000000000000",23588 => "0000000000000000",
23589 => "0000000000000000",23590 => "0000000000000000",
23591 => "0000000000000000",23592 => "0000000000000000",
23593 => "0000000000000000",23594 => "0000000000000000",
23595 => "0000000000000000",23596 => "0000000000000000",
23597 => "0000000000000000",23598 => "0000000000000000",
23599 => "0000000000000000",23600 => "0000000000000000",
23601 => "0000000000000000",23602 => "0000000000000000",
23603 => "0000000000000000",23604 => "0000000000000000",
23605 => "0000000000000000",23606 => "0000000000000000",
23607 => "0000000000000000",23608 => "0000000000000000",
23609 => "0000000000000000",23610 => "0000000000000000",
23611 => "0000000000000000",23612 => "0000000000000000",
23613 => "0000000000000000",23614 => "0000000000000000",
23615 => "0000000000000000",23616 => "0000000000000000",
23617 => "0000000000000000",23618 => "0000000000000000",
23619 => "0000000000000000",23620 => "0000000000000000",
23621 => "0000000000000000",23622 => "0000000000000000",
23623 => "0000000000000000",23624 => "0000000000000000",
23625 => "0000000000000000",23626 => "0000000000000000",
23627 => "0000000000000000",23628 => "0000000000000000",
23629 => "0000000000000000",23630 => "0000000000000000",
23631 => "0000000000000000",23632 => "0000000000000000",
23633 => "0000000000000000",23634 => "0000000000000000",
23635 => "0000000000000000",23636 => "0000000000000000",
23637 => "0000000000000000",23638 => "0000000000000000",
23639 => "0000000000000000",23640 => "0000000000000000",
23641 => "0000000000000000",23642 => "0000000000000000",
23643 => "0000000000000000",23644 => "0000000000000000",
23645 => "0000000000000000",23646 => "0000000000000000",
23647 => "0000000000000000",23648 => "0000000000000000",
23649 => "0000000000000000",23650 => "0000000000000000",
23651 => "0000000000000000",23652 => "0000000000000000",
23653 => "0000000000000000",23654 => "0000000000000000",
23655 => "0000000000000000",23656 => "0000000000000000",
23657 => "0000000000000000",23658 => "0000000000000000",
23659 => "0000000000000000",23660 => "0000000000000000",
23661 => "0000000000000000",23662 => "0000000000000000",
23663 => "0000000000000000",23664 => "0000000000000000",
23665 => "0000000000000000",23666 => "0000000000000000",
23667 => "0000000000000000",23668 => "0000000000000000",
23669 => "0000000000000000",23670 => "0000000000000000",
23671 => "0000000000000000",23672 => "0000000000000000",
23673 => "0000000000000000",23674 => "0000000000000000",
23675 => "0000000000000000",23676 => "0000000000000000",
23677 => "0000000000000000",23678 => "0000000000000000",
23679 => "0000000000000000",23680 => "0000000000000000",
23681 => "0000000000000000",23682 => "0000000000000000",
23683 => "0000000000000000",23684 => "0000000000000000",
23685 => "0000000000000000",23686 => "0000000000000000",
23687 => "0000000000000000",23688 => "0000000000000000",
23689 => "0000000000000000",23690 => "0000000000000000",
23691 => "0000000000000000",23692 => "0000000000000000",
23693 => "0000000000000000",23694 => "0000000000000000",
23695 => "0000000000000000",23696 => "0000000000000000",
23697 => "0000000000000000",23698 => "0000000000000000",
23699 => "0000000000000000",23700 => "0000000000000000",
23701 => "0000000000000000",23702 => "0000000000000000",
23703 => "0000000000000000",23704 => "0000000000000000",
23705 => "0000000000000000",23706 => "0000000000000000",
23707 => "0000000000000000",23708 => "0000000000000000",
23709 => "0000000000000000",23710 => "0000000000000000",
23711 => "0000000000000000",23712 => "0000000000000000",
23713 => "0000000000000000",23714 => "0000000000000000",
23715 => "0000000000000000",23716 => "0000000000000000",
23717 => "0000000000000000",23718 => "0000000000000000",
23719 => "0000000000000000",23720 => "0000000000000000",
23721 => "0000000000000000",23722 => "0000000000000000",
23723 => "0000000000000000",23724 => "0000000000000000",
23725 => "0000000000000000",23726 => "0000000000000000",
23727 => "0000000000000000",23728 => "0000000000000000",
23729 => "0000000000000000",23730 => "0000000000000000",
23731 => "0000000000000000",23732 => "0000000000000000",
23733 => "0000000000000000",23734 => "0000000000000000",
23735 => "0000000000000000",23736 => "0000000000000000",
23737 => "0000000000000000",23738 => "0000000000000000",
23739 => "0000000000000000",23740 => "0000000000000000",
23741 => "0000000000000000",23742 => "0000000000000000",
23743 => "0000000000000000",23744 => "0000000000000000",
23745 => "0000000000000000",23746 => "0000000000000000",
23747 => "0000000000000000",23748 => "0000000000000000",
23749 => "0000000000000000",23750 => "0000000000000000",
23751 => "0000000000000000",23752 => "0000000000000000",
23753 => "0000000000000000",23754 => "0000000000000000",
23755 => "0000000000000000",23756 => "0000000000000000",
23757 => "0000000000000000",23758 => "0000000000000000",
23759 => "0000000000000000",23760 => "0000000000000000",
23761 => "0000000000000000",23762 => "0000000000000000",
23763 => "0000000000000000",23764 => "0000000000000000",
23765 => "0000000000000000",23766 => "0000000000000000",
23767 => "0000000000000000",23768 => "0000000000000000",
23769 => "0000000000000000",23770 => "0000000000000000",
23771 => "0000000000000000",23772 => "0000000000000000",
23773 => "0000000000000000",23774 => "0000000000000000",
23775 => "0000000000000000",23776 => "0000000000000000",
23777 => "0000000000000000",23778 => "0000000000000000",
23779 => "0000000000000000",23780 => "0000000000000000",
23781 => "0000000000000000",23782 => "0000000000000000",
23783 => "0000000000000000",23784 => "0000000000000000",
23785 => "0000000000000000",23786 => "0000000000000000",
23787 => "0000000000000000",23788 => "0000000000000000",
23789 => "0000000000000000",23790 => "0000000000000000",
23791 => "0000000000000000",23792 => "0000000000000000",
23793 => "0000000000000000",23794 => "0000000000000000",
23795 => "0000000000000000",23796 => "0000000000000000",
23797 => "0000000000000000",23798 => "0000000000000000",
23799 => "0000000000000000",23800 => "0000000000000000",
23801 => "0000000000000000",23802 => "0000000000000000",
23803 => "0000000000000000",23804 => "0000000000000000",
23805 => "0000000000000000",23806 => "0000000000000000",
23807 => "0000000000000000",23808 => "0000000000000000",
23809 => "0000000000000000",23810 => "0000000000000000",
23811 => "0000000000000000",23812 => "0000000000000000",
23813 => "0000000000000000",23814 => "0000000000000000",
23815 => "0000000000000000",23816 => "0000000000000000",
23817 => "0000000000000000",23818 => "0000000000000000",
23819 => "0000000000000000",23820 => "0000000000000000",
23821 => "0000000000000000",23822 => "0000000000000000",
23823 => "0000000000000000",23824 => "0000000000000000",
23825 => "0000000000000000",23826 => "0000000000000000",
23827 => "0000000000000000",23828 => "0000000000000000",
23829 => "0000000000000000",23830 => "0000000000000000",
23831 => "0000000000000000",23832 => "0000000000000000",
23833 => "0000000000000000",23834 => "0000000000000000",
23835 => "0000000000000000",23836 => "0000000000000000",
23837 => "0000000000000000",23838 => "0000000000000000",
23839 => "0000000000000000",23840 => "0000000000000000",
23841 => "0000000000000000",23842 => "0000000000000000",
23843 => "0000000000000000",23844 => "0000000000000000",
23845 => "0000000000000000",23846 => "0000000000000000",
23847 => "0000000000000000",23848 => "0000000000000000",
23849 => "0000000000000000",23850 => "0000000000000000",
23851 => "0000000000000000",23852 => "0000000000000000",
23853 => "0000000000000000",23854 => "0000000000000000",
23855 => "0000000000000000",23856 => "0000000000000000",
23857 => "0000000000000000",23858 => "0000000000000000",
23859 => "0000000000000000",23860 => "0000000000000000",
23861 => "0000000000000000",23862 => "0000000000000000",
23863 => "0000000000000000",23864 => "0000000000000000",
23865 => "0000000000000000",23866 => "0000000000000000",
23867 => "0000000000000000",23868 => "0000000000000000",
23869 => "0000000000000000",23870 => "0000000000000000",
23871 => "0000000000000000",23872 => "0000000000000000",
23873 => "0000000000000000",23874 => "0000000000000000",
23875 => "0000000000000000",23876 => "0000000000000000",
23877 => "0000000000000000",23878 => "0000000000000000",
23879 => "0000000000000000",23880 => "0000000000000000",
23881 => "0000000000000000",23882 => "0000000000000000",
23883 => "0000000000000000",23884 => "0000000000000000",
23885 => "0000000000000000",23886 => "0000000000000000",
23887 => "0000000000000000",23888 => "0000000000000000",
23889 => "0000000000000000",23890 => "0000000000000000",
23891 => "0000000000000000",23892 => "0000000000000000",
23893 => "0000000000000000",23894 => "0000000000000000",
23895 => "0000000000000000",23896 => "0000000000000000",
23897 => "0000000000000000",23898 => "0000000000000000",
23899 => "0000000000000000",23900 => "0000000000000000",
23901 => "0000000000000000",23902 => "0000000000000000",
23903 => "0000000000000000",23904 => "0000000000000000",
23905 => "0000000000000000",23906 => "0000000000000000",
23907 => "0000000000000000",23908 => "0000000000000000",
23909 => "0000000000000000",23910 => "0000000000000000",
23911 => "0000000000000000",23912 => "0000000000000000",
23913 => "0000000000000000",23914 => "0000000000000000",
23915 => "0000000000000000",23916 => "0000000000000000",
23917 => "0000000000000000",23918 => "0000000000000000",
23919 => "0000000000000000",23920 => "0000000000000000",
23921 => "0000000000000000",23922 => "0000000000000000",
23923 => "0000000000000000",23924 => "0000000000000000",
23925 => "0000000000000000",23926 => "0000000000000000",
23927 => "0000000000000000",23928 => "0000000000000000",
23929 => "0000000000000000",23930 => "0000000000000000",
23931 => "0000000000000000",23932 => "0000000000000000",
23933 => "0000000000000000",23934 => "0000000000000000",
23935 => "0000000000000000",23936 => "0000000000000000",
23937 => "0000000000000000",23938 => "0000000000000000",
23939 => "0000000000000000",23940 => "0000000000000000",
23941 => "0000000000000000",23942 => "0000000000000000",
23943 => "0000000000000000",23944 => "0000000000000000",
23945 => "0000000000000000",23946 => "0000000000000000",
23947 => "0000000000000000",23948 => "0000000000000000",
23949 => "0000000000000000",23950 => "0000000000000000",
23951 => "0000000000000000",23952 => "0000000000000000",
23953 => "0000000000000000",23954 => "0000000000000000",
23955 => "0000000000000000",23956 => "0000000000000000",
23957 => "0000000000000000",23958 => "0000000000000000",
23959 => "0000000000000000",23960 => "0000000000000000",
23961 => "0000000000000000",23962 => "0000000000000000",
23963 => "0000000000000000",23964 => "0000000000000000",
23965 => "0000000000000000",23966 => "0000000000000000",
23967 => "0000000000000000",23968 => "0000000000000000",
23969 => "0000000000000000",23970 => "0000000000000000",
23971 => "0000000000000000",23972 => "0000000000000000",
23973 => "0000000000000000",23974 => "0000000000000000",
23975 => "0000000000000000",23976 => "0000000000000000",
23977 => "0000000000000000",23978 => "0000000000000000",
23979 => "0000000000000000",23980 => "0000000000000000",
23981 => "0000000000000000",23982 => "0000000000000000",
23983 => "0000000000000000",23984 => "0000000000000000",
23985 => "0000000000000000",23986 => "0000000000000000",
23987 => "0000000000000000",23988 => "0000000000000000",
23989 => "0000000000000000",23990 => "0000000000000000",
23991 => "0000000000000000",23992 => "0000000000000000",
23993 => "0000000000000000",23994 => "0000000000000000",
23995 => "0000000000000000",23996 => "0000000000000000",
23997 => "0000000000000000",23998 => "0000000000000000",
23999 => "0000000000000000",24000 => "0000000000000000",
24001 => "0000000000000000",24002 => "0000000000000000",
24003 => "0000000000000000",24004 => "0000000000000000",
24005 => "0000000000000000",24006 => "0000000000000000",
24007 => "0000000000000000",24008 => "0000000000000000",
24009 => "0000000000000000",24010 => "0000000000000000",
24011 => "0000000000000000",24012 => "0000000000000000",
24013 => "0000000000000000",24014 => "0000000000000000",
24015 => "0000000000000000",24016 => "0000000000000000",
24017 => "0000000000000000",24018 => "0000000000000000",
24019 => "0000000000000000",24020 => "0000000000000000",
24021 => "0000000000000000",24022 => "0000000000000000",
24023 => "0000000000000000",24024 => "0000000000000000",
24025 => "0000000000000000",24026 => "0000000000000000",
24027 => "0000000000000000",24028 => "0000000000000000",
24029 => "0000000000000000",24030 => "0000000000000000",
24031 => "0000000000000000",24032 => "0000000000000000",
24033 => "0000000000000000",24034 => "0000000000000000",
24035 => "0000000000000000",24036 => "0000000000000000",
24037 => "0000000000000000",24038 => "0000000000000000",
24039 => "0000000000000000",24040 => "0000000000000000",
24041 => "0000000000000000",24042 => "0000000000000000",
24043 => "0000000000000000",24044 => "0000000000000000",
24045 => "0000000000000000",24046 => "0000000000000000",
24047 => "0000000000000000",24048 => "0000000000000000",
24049 => "0000000000000000",24050 => "0000000000000000",
24051 => "0000000000000000",24052 => "0000000000000000",
24053 => "0000000000000000",24054 => "0000000000000000",
24055 => "0000000000000000",24056 => "0000000000000000",
24057 => "0000000000000000",24058 => "0000000000000000",
24059 => "0000000000000000",24060 => "0000000000000000",
24061 => "0000000000000000",24062 => "0000000000000000",
24063 => "0000000000000000",24064 => "0000000000000000",
24065 => "0000000000000000",24066 => "0000000000000000",
24067 => "0000000000000000",24068 => "0000000000000000",
24069 => "0000000000000000",24070 => "0000000000000000",
24071 => "0000000000000000",24072 => "0000000000000000",
24073 => "0000000000000000",24074 => "0000000000000000",
24075 => "0000000000000000",24076 => "0000000000000000",
24077 => "0000000000000000",24078 => "0000000000000000",
24079 => "0000000000000000",24080 => "0000000000000000",
24081 => "0000000000000000",24082 => "0000000000000000",
24083 => "0000000000000000",24084 => "0000000000000000",
24085 => "0000000000000000",24086 => "0000000000000000",
24087 => "0000000000000000",24088 => "0000000000000000",
24089 => "0000000000000000",24090 => "0000000000000000",
24091 => "0000000000000000",24092 => "0000000000000000",
24093 => "0000000000000000",24094 => "0000000000000000",
24095 => "0000000000000000",24096 => "0000000000000000",
24097 => "0000000000000000",24098 => "0000000000000000",
24099 => "0000000000000000",24100 => "0000000000000000",
24101 => "0000000000000000",24102 => "0000000000000000",
24103 => "0000000000000000",24104 => "0000000000000000",
24105 => "0000000000000000",24106 => "0000000000000000",
24107 => "0000000000000000",24108 => "0000000000000000",
24109 => "0000000000000000",24110 => "0000000000000000",
24111 => "0000000000000000",24112 => "0000000000000000",
24113 => "0000000000000000",24114 => "0000000000000000",
24115 => "0000000000000000",24116 => "0000000000000000",
24117 => "0000000000000000",24118 => "0000000000000000",
24119 => "0000000000000000",24120 => "0000000000000000",
24121 => "0000000000000000",24122 => "0000000000000000",
24123 => "0000000000000000",24124 => "0000000000000000",
24125 => "0000000000000000",24126 => "0000000000000000",
24127 => "0000000000000000",24128 => "0000000000000000",
24129 => "0000000000000000",24130 => "0000000000000000",
24131 => "0000000000000000",24132 => "0000000000000000",
24133 => "0000000000000000",24134 => "0000000000000000",
24135 => "0000000000000000",24136 => "0000000000000000",
24137 => "0000000000000000",24138 => "0000000000000000",
24139 => "0000000000000000",24140 => "0000000000000000",
24141 => "0000000000000000",24142 => "0000000000000000",
24143 => "0000000000000000",24144 => "0000000000000000",
24145 => "0000000000000000",24146 => "0000000000000000",
24147 => "0000000000000000",24148 => "0000000000000000",
24149 => "0000000000000000",24150 => "0000000000000000",
24151 => "0000000000000000",24152 => "0000000000000000",
24153 => "0000000000000000",24154 => "0000000000000000",
24155 => "0000000000000000",24156 => "0000000000000000",
24157 => "0000000000000000",24158 => "0000000000000000",
24159 => "0000000000000000",24160 => "0000000000000000",
24161 => "0000000000000000",24162 => "0000000000000000",
24163 => "0000000000000000",24164 => "0000000000000000",
24165 => "0000000000000000",24166 => "0000000000000000",
24167 => "0000000000000000",24168 => "0000000000000000",
24169 => "0000000000000000",24170 => "0000000000000000",
24171 => "0000000000000000",24172 => "0000000000000000",
24173 => "0000000000000000",24174 => "0000000000000000",
24175 => "0000000000000000",24176 => "0000000000000000",
24177 => "0000000000000000",24178 => "0000000000000000",
24179 => "0000000000000000",24180 => "0000000000000000",
24181 => "0000000000000000",24182 => "0000000000000000",
24183 => "0000000000000000",24184 => "0000000000000000",
24185 => "0000000000000000",24186 => "0000000000000000",
24187 => "0000000000000000",24188 => "0000000000000000",
24189 => "0000000000000000",24190 => "0000000000000000",
24191 => "0000000000000000",24192 => "0000000000000000",
24193 => "0000000000000000",24194 => "0000000000000000",
24195 => "0000000000000000",24196 => "0000000000000000",
24197 => "0000000000000000",24198 => "0000000000000000",
24199 => "0000000000000000",24200 => "0000000000000000",
24201 => "0000000000000000",24202 => "0000000000000000",
24203 => "0000000000000000",24204 => "0000000000000000",
24205 => "0000000000000000",24206 => "0000000000000000",
24207 => "0000000000000000",24208 => "0000000000000000",
24209 => "0000000000000000",24210 => "0000000000000000",
24211 => "0000000000000000",24212 => "0000000000000000",
24213 => "0000000000000000",24214 => "0000000000000000",
24215 => "0000000000000000",24216 => "0000000000000000",
24217 => "0000000000000000",24218 => "0000000000000000",
24219 => "0000000000000000",24220 => "0000000000000000",
24221 => "0000000000000000",24222 => "0000000000000000",
24223 => "0000000000000000",24224 => "0000000000000000",
24225 => "0000000000000000",24226 => "0000000000000000",
24227 => "0000000000000000",24228 => "0000000000000000",
24229 => "0000000000000000",24230 => "0000000000000000",
24231 => "0000000000000000",24232 => "0000000000000000",
24233 => "0000000000000000",24234 => "0000000000000000",
24235 => "0000000000000000",24236 => "0000000000000000",
24237 => "0000000000000000",24238 => "0000000000000000",
24239 => "0000000000000000",24240 => "0000000000000000",
24241 => "0000000000000000",24242 => "0000000000000000",
24243 => "0000000000000000",24244 => "0000000000000000",
24245 => "0000000000000000",24246 => "0000000000000000",
24247 => "0000000000000000",24248 => "0000000000000000",
24249 => "0000000000000000",24250 => "0000000000000000",
24251 => "0000000000000000",24252 => "0000000000000000",
24253 => "0000000000000000",24254 => "0000000000000000",
24255 => "0000000000000000",24256 => "0000000000000000",
24257 => "0000000000000000",24258 => "0000000000000000",
24259 => "0000000000000000",24260 => "0000000000000000",
24261 => "0000000000000000",24262 => "0000000000000000",
24263 => "0000000000000000",24264 => "0000000000000000",
24265 => "0000000000000000",24266 => "0000000000000000",
24267 => "0000000000000000",24268 => "0000000000000000",
24269 => "0000000000000000",24270 => "0000000000000000",
24271 => "0000000000000000",24272 => "0000000000000000",
24273 => "0000000000000000",24274 => "0000000000000000",
24275 => "0000000000000000",24276 => "0000000000000000",
24277 => "0000000000000000",24278 => "0000000000000000",
24279 => "0000000000000000",24280 => "0000000000000000",
24281 => "0000000000000000",24282 => "0000000000000000",
24283 => "0000000000000000",24284 => "0000000000000000",
24285 => "0000000000000000",24286 => "0000000000000000",
24287 => "0000000000000000",24288 => "0000000000000000",
24289 => "0000000000000000",24290 => "0000000000000000",
24291 => "0000000000000000",24292 => "0000000000000000",
24293 => "0000000000000000",24294 => "0000000000000000",
24295 => "0000000000000000",24296 => "0000000000000000",
24297 => "0000000000000000",24298 => "0000000000000000",
24299 => "0000000000000000",24300 => "0000000000000000",
24301 => "0000000000000000",24302 => "0000000000000000",
24303 => "0000000000000000",24304 => "0000000000000000",
24305 => "0000000000000000",24306 => "0000000000000000",
24307 => "0000000000000000",24308 => "0000000000000000",
24309 => "0000000000000000",24310 => "0000000000000000",
24311 => "0000000000000000",24312 => "0000000000000000",
24313 => "0000000000000000",24314 => "0000000000000000",
24315 => "0000000000000000",24316 => "0000000000000000",
24317 => "0000000000000000",24318 => "0000000000000000",
24319 => "0000000000000000",24320 => "0000000000000000",
24321 => "0000000000000000",24322 => "0000000000000000",
24323 => "0000000000000000",24324 => "0000000000000000",
24325 => "0000000000000000",24326 => "0000000000000000",
24327 => "0000000000000000",24328 => "0000000000000000",
24329 => "0000000000000000",24330 => "0000000000000000",
24331 => "0000000000000000",24332 => "0000000000000000",
24333 => "0000000000000000",24334 => "0000000000000000",
24335 => "0000000000000000",24336 => "0000000000000000",
24337 => "0000000000000000",24338 => "0000000000000000",
24339 => "0000000000000000",24340 => "0000000000000000",
24341 => "0000000000000000",24342 => "0000000000000000",
24343 => "0000000000000000",24344 => "0000000000000000",
24345 => "0000000000000000",24346 => "0000000000000000",
24347 => "0000000000000000",24348 => "0000000000000000",
24349 => "0000000000000000",24350 => "0000000000000000",
24351 => "0000000000000000",24352 => "0000000000000000",
24353 => "0000000000000000",24354 => "0000000000000000",
24355 => "0000000000000000",24356 => "0000000000000000",
24357 => "0000000000000000",24358 => "0000000000000000",
24359 => "0000000000000000",24360 => "0000000000000000",
24361 => "0000000000000000",24362 => "0000000000000000",
24363 => "0000000000000000",24364 => "0000000000000000",
24365 => "0000000000000000",24366 => "0000000000000000",
24367 => "0000000000000000",24368 => "0000000000000000",
24369 => "0000000000000000",24370 => "0000000000000000",
24371 => "0000000000000000",24372 => "0000000000000000",
24373 => "0000000000000000",24374 => "0000000000000000",
24375 => "0000000000000000",24376 => "0000000000000000",
24377 => "0000000000000000",24378 => "0000000000000000",
24379 => "0000000000000000",24380 => "0000000000000000",
24381 => "0000000000000000",24382 => "0000000000000000",
24383 => "0000000000000000",24384 => "0000000000000000",
24385 => "0000000000000000",24386 => "0000000000000000",
24387 => "0000000000000000",24388 => "0000000000000000",
24389 => "0000000000000000",24390 => "0000000000000000",
24391 => "0000000000000000",24392 => "0000000000000000",
24393 => "0000000000000000",24394 => "0000000000000000",
24395 => "0000000000000000",24396 => "0000000000000000",
24397 => "0000000000000000",24398 => "0000000000000000",
24399 => "0000000000000000",24400 => "0000000000000000",
24401 => "0000000000000000",24402 => "0000000000000000",
24403 => "0000000000000000",24404 => "0000000000000000",
24405 => "0000000000000000",24406 => "0000000000000000",
24407 => "0000000000000000",24408 => "0000000000000000",
24409 => "0000000000000000",24410 => "0000000000000000",
24411 => "0000000000000000",24412 => "0000000000000000",
24413 => "0000000000000000",24414 => "0000000000000000",
24415 => "0000000000000000",24416 => "0000000000000000",
24417 => "0000000000000000",24418 => "0000000000000000",
24419 => "0000000000000000",24420 => "0000000000000000",
24421 => "0000000000000000",24422 => "0000000000000000",
24423 => "0000000000000000",24424 => "0000000000000000",
24425 => "0000000000000000",24426 => "0000000000000000",
24427 => "0000000000000000",24428 => "0000000000000000",
24429 => "0000000000000000",24430 => "0000000000000000",
24431 => "0000000000000000",24432 => "0000000000000000",
24433 => "0000000000000000",24434 => "0000000000000000",
24435 => "0000000000000000",24436 => "0000000000000000",
24437 => "0000000000000000",24438 => "0000000000000000",
24439 => "0000000000000000",24440 => "0000000000000000",
24441 => "0000000000000000",24442 => "0000000000000000",
24443 => "0000000000000000",24444 => "0000000000000000",
24445 => "0000000000000000",24446 => "0000000000000000",
24447 => "0000000000000000",24448 => "0000000000000000",
24449 => "0000000000000000",24450 => "0000000000000000",
24451 => "0000000000000000",24452 => "0000000000000000",
24453 => "0000000000000000",24454 => "0000000000000000",
24455 => "0000000000000000",24456 => "0000000000000000",
24457 => "0000000000000000",24458 => "0000000000000000",
24459 => "0000000000000000",24460 => "0000000000000000",
24461 => "0000000000000000",24462 => "0000000000000000",
24463 => "0000000000000000",24464 => "0000000000000000",
24465 => "0000000000000000",24466 => "0000000000000000",
24467 => "0000000000000000",24468 => "0000000000000000",
24469 => "0000000000000000",24470 => "0000000000000000",
24471 => "0000000000000000",24472 => "0000000000000000",
24473 => "0000000000000000",24474 => "0000000000000000",
24475 => "0000000000000000",24476 => "0000000000000000",
24477 => "0000000000000000",24478 => "0000000000000000",
24479 => "0000000000000000",24480 => "0000000000000000",
24481 => "0000000000000000",24482 => "0000000000000000",
24483 => "0000000000000000",24484 => "0000000000000000",
24485 => "0000000000000000",24486 => "0000000000000000",
24487 => "0000000000000000",24488 => "0000000000000000",
24489 => "0000000000000000",24490 => "0000000000000000",
24491 => "0000000000000000",24492 => "0000000000000000",
24493 => "0000000000000000",24494 => "0000000000000000",
24495 => "0000000000000000",24496 => "0000000000000000",
24497 => "0000000000000000",24498 => "0000000000000000",
24499 => "0000000000000000",24500 => "0000000000000000",
24501 => "0000000000000000",24502 => "0000000000000000",
24503 => "0000000000000000",24504 => "0000000000000000",
24505 => "0000000000000000",24506 => "0000000000000000",
24507 => "0000000000000000",24508 => "0000000000000000",
24509 => "0000000000000000",24510 => "0000000000000000",
24511 => "0000000000000000",24512 => "0000000000000000",
24513 => "0000000000000000",24514 => "0000000000000000",
24515 => "0000000000000000",24516 => "0000000000000000",
24517 => "0000000000000000",24518 => "0000000000000000",
24519 => "0000000000000000",24520 => "0000000000000000",
24521 => "0000000000000000",24522 => "0000000000000000",
24523 => "0000000000000000",24524 => "0000000000000000",
24525 => "0000000000000000",24526 => "0000000000000000",
24527 => "0000000000000000",24528 => "0000000000000000",
24529 => "0000000000000000",24530 => "0000000000000000",
24531 => "0000000000000000",24532 => "0000000000000000",
24533 => "0000000000000000",24534 => "0000000000000000",
24535 => "0000000000000000",24536 => "0000000000000000",
24537 => "0000000000000000",24538 => "0000000000000000",
24539 => "0000000000000000",24540 => "0000000000000000",
24541 => "0000000000000000",24542 => "0000000000000000",
24543 => "0000000000000000",24544 => "0000000000000000",
24545 => "0000000000000000",24546 => "0000000000000000",
24547 => "0000000000000000",24548 => "0000000000000000",
24549 => "0000000000000000",24550 => "0000000000000000",
24551 => "0000000000000000",24552 => "0000000000000000",
24553 => "0000000000000000",24554 => "0000000000000000",
24555 => "0000000000000000",24556 => "0000000000000000",
24557 => "0000000000000000",24558 => "0000000000000000",
24559 => "0000000000000000",24560 => "0000000000000000",
24561 => "0000000000000000",24562 => "0000000000000000",
24563 => "0000000000000000",24564 => "0000000000000000",
24565 => "0000000000000000",24566 => "0000000000000000",
24567 => "0000000000000000",24568 => "0000000000000000",
24569 => "0000000000000000",24570 => "0000000000000000",
24571 => "0000000000000000",24572 => "0000000000000000",
24573 => "0000000000000000",24574 => "0000000000000000",
24575 => "0000000000000000",24576 => "0000000000000000",
24577 => "0000000000000000",24578 => "0000000000000000",
24579 => "0000000000000000",24580 => "0000000000000000",
24581 => "0000000000000000",24582 => "0000000000000000",
24583 => "0000000000000000",24584 => "0000000000000000",
24585 => "0000000000000000",24586 => "0000000000000000",
24587 => "0000000000000000",24588 => "0000000000000000",
24589 => "0000000000000000",24590 => "0000000000000000",
24591 => "0000000000000000",24592 => "0000000000000000",
24593 => "0000000000000000",24594 => "0000000000000000",
24595 => "0000000000000000",24596 => "0000000000000000",
24597 => "0000000000000000",24598 => "0000000000000000",
24599 => "0000000000000000",24600 => "0000000000000000",
24601 => "0000000000000000",24602 => "0000000000000000",
24603 => "0000000000000000",24604 => "0000000000000000",
24605 => "0000000000000000",24606 => "0000000000000000",
24607 => "0000000000000000",24608 => "0000000000000000",
24609 => "0000000000000000",24610 => "0000000000000000",
24611 => "0000000000000000",24612 => "0000000000000000",
24613 => "0000000000000000",24614 => "0000000000000000",
24615 => "0000000000000000",24616 => "0000000000000000",
24617 => "0000000000000000",24618 => "0000000000000000",
24619 => "0000000000000000",24620 => "0000000000000000",
24621 => "0000000000000000",24622 => "0000000000000000",
24623 => "0000000000000000",24624 => "0000000000000000",
24625 => "0000000000000000",24626 => "0000000000000000",
24627 => "0000000000000000",24628 => "0000000000000000",
24629 => "0000000000000000",24630 => "0000000000000000",
24631 => "0000000000000000",24632 => "0000000000000000",
24633 => "0000000000000000",24634 => "0000000000000000",
24635 => "0000000000000000",24636 => "0000000000000000",
24637 => "0000000000000000",24638 => "0000000000000000",
24639 => "0000000000000000",24640 => "0000000000000000",
24641 => "0000000000000000",24642 => "0000000000000000",
24643 => "0000000000000000",24644 => "0000000000000000",
24645 => "0000000000000000",24646 => "0000000000000000",
24647 => "0000000000000000",24648 => "0000000000000000",
24649 => "0000000000000000",24650 => "0000000000000000",
24651 => "0000000000000000",24652 => "0000000000000000",
24653 => "0000000000000000",24654 => "0000000000000000",
24655 => "0000000000000000",24656 => "0000000000000000",
24657 => "0000000000000000",24658 => "0000000000000000",
24659 => "0000000000000000",24660 => "0000000000000000",
24661 => "0000000000000000",24662 => "0000000000000000",
24663 => "0000000000000000",24664 => "0000000000000000",
24665 => "0000000000000000",24666 => "0000000000000000",
24667 => "0000000000000000",24668 => "0000000000000000",
24669 => "0000000000000000",24670 => "0000000000000000",
24671 => "0000000000000000",24672 => "0000000000000000",
24673 => "0000000000000000",24674 => "0000000000000000",
24675 => "0000000000000000",24676 => "0000000000000000",
24677 => "0000000000000000",24678 => "0000000000000000",
24679 => "0000000000000000",24680 => "0000000000000000",
24681 => "0000000000000000",24682 => "0000000000000000",
24683 => "0000000000000000",24684 => "0000000000000000",
24685 => "0000000000000000",24686 => "0000000000000000",
24687 => "0000000000000000",24688 => "0000000000000000",
24689 => "0000000000000000",24690 => "0000000000000000",
24691 => "0000000000000000",24692 => "0000000000000000",
24693 => "0000000000000000",24694 => "0000000000000000",
24695 => "0000000000000000",24696 => "0000000000000000",
24697 => "0000000000000000",24698 => "0000000000000000",
24699 => "0000000000000000",24700 => "0000000000000000",
24701 => "0000000000000000",24702 => "0000000000000000",
24703 => "0000000000000000",24704 => "0000000000000000",
24705 => "0000000000000000",24706 => "0000000000000000",
24707 => "0000000000000000",24708 => "0000000000000000",
24709 => "0000000000000000",24710 => "0000000000000000",
24711 => "0000000000000000",24712 => "0000000000000000",
24713 => "0000000000000000",24714 => "0000000000000000",
24715 => "0000000000000000",24716 => "0000000000000000",
24717 => "0000000000000000",24718 => "0000000000000000",
24719 => "0000000000000000",24720 => "0000000000000000",
24721 => "0000000000000000",24722 => "0000000000000000",
24723 => "0000000000000000",24724 => "0000000000000000",
24725 => "0000000000000000",24726 => "0000000000000000",
24727 => "0000000000000000",24728 => "0000000000000000",
24729 => "0000000000000000",24730 => "0000000000000000",
24731 => "0000000000000000",24732 => "0000000000000000",
24733 => "0000000000000000",24734 => "0000000000000000",
24735 => "0000000000000000",24736 => "0000000000000000",
24737 => "0000000000000000",24738 => "0000000000000000",
24739 => "0000000000000000",24740 => "0000000000000000",
24741 => "0000000000000000",24742 => "0000000000000000",
24743 => "0000000000000000",24744 => "0000000000000000",
24745 => "0000000000000000",24746 => "0000000000000000",
24747 => "0000000000000000",24748 => "0000000000000000",
24749 => "0000000000000000",24750 => "0000000000000000",
24751 => "0000000000000000",24752 => "0000000000000000",
24753 => "0000000000000000",24754 => "0000000000000000",
24755 => "0000000000000000",24756 => "0000000000000000",
24757 => "0000000000000000",24758 => "0000000000000000",
24759 => "0000000000000000",24760 => "0000000000000000",
24761 => "0000000000000000",24762 => "0000000000000000",
24763 => "0000000000000000",24764 => "0000000000000000",
24765 => "0000000000000000",24766 => "0000000000000000",
24767 => "0000000000000000",24768 => "0000000000000000",
24769 => "0000000000000000",24770 => "0000000000000000",
24771 => "0000000000000000",24772 => "0000000000000000",
24773 => "0000000000000000",24774 => "0000000000000000",
24775 => "0000000000000000",24776 => "0000000000000000",
24777 => "0000000000000000",24778 => "0000000000000000",
24779 => "0000000000000000",24780 => "0000000000000000",
24781 => "0000000000000000",24782 => "0000000000000000",
24783 => "0000000000000000",24784 => "0000000000000000",
24785 => "0000000000000000",24786 => "0000000000000000",
24787 => "0000000000000000",24788 => "0000000000000000",
24789 => "0000000000000000",24790 => "0000000000000000",
24791 => "0000000000000000",24792 => "0000000000000000",
24793 => "0000000000000000",24794 => "0000000000000000",
24795 => "0000000000000000",24796 => "0000000000000000",
24797 => "0000000000000000",24798 => "0000000000000000",
24799 => "0000000000000000",24800 => "0000000000000000",
24801 => "0000000000000000",24802 => "0000000000000000",
24803 => "0000000000000000",24804 => "0000000000000000",
24805 => "0000000000000000",24806 => "0000000000000000",
24807 => "0000000000000000",24808 => "0000000000000000",
24809 => "0000000000000000",24810 => "0000000000000000",
24811 => "0000000000000000",24812 => "0000000000000000",
24813 => "0000000000000000",24814 => "0000000000000000",
24815 => "0000000000000000",24816 => "0000000000000000",
24817 => "0000000000000000",24818 => "0000000000000000",
24819 => "0000000000000000",24820 => "0000000000000000",
24821 => "0000000000000000",24822 => "0000000000000000",
24823 => "0000000000000000",24824 => "0000000000000000",
24825 => "0000000000000000",24826 => "0000000000000000",
24827 => "0000000000000000",24828 => "0000000000000000",
24829 => "0000000000000000",24830 => "0000000000000000",
24831 => "0000000000000000",24832 => "0000000000000000",
24833 => "0000000000000000",24834 => "0000000000000000",
24835 => "0000000000000000",24836 => "0000000000000000",
24837 => "0000000000000000",24838 => "0000000000000000",
24839 => "0000000000000000",24840 => "0000000000000000",
24841 => "0000000000000000",24842 => "0000000000000000",
24843 => "0000000000000000",24844 => "0000000000000000",
24845 => "0000000000000000",24846 => "0000000000000000",
24847 => "0000000000000000",24848 => "0000000000000000",
24849 => "0000000000000000",24850 => "0000000000000000",
24851 => "0000000000000000",24852 => "0000000000000000",
24853 => "0000000000000000",24854 => "0000000000000000",
24855 => "0000000000000000",24856 => "0000000000000000",
24857 => "0000000000000000",24858 => "0000000000000000",
24859 => "0000000000000000",24860 => "0000000000000000",
24861 => "0000000000000000",24862 => "0000000000000000",
24863 => "0000000000000000",24864 => "0000000000000000",
24865 => "0000000000000000",24866 => "0000000000000000",
24867 => "0000000000000000",24868 => "0000000000000000",
24869 => "0000000000000000",24870 => "0000000000000000",
24871 => "0000000000000000",24872 => "0000000000000000",
24873 => "0000000000000000",24874 => "0000000000000000",
24875 => "0000000000000000",24876 => "0000000000000000",
24877 => "0000000000000000",24878 => "0000000000000000",
24879 => "0000000000000000",24880 => "0000000000000000",
24881 => "0000000000000000",24882 => "0000000000000000",
24883 => "0000000000000000",24884 => "0000000000000000",
24885 => "0000000000000000",24886 => "0000000000000000",
24887 => "0000000000000000",24888 => "0000000000000000",
24889 => "0000000000000000",24890 => "0000000000000000",
24891 => "0000000000000000",24892 => "0000000000000000",
24893 => "0000000000000000",24894 => "0000000000000000",
24895 => "0000000000000000",24896 => "0000000000000000",
24897 => "0000000000000000",24898 => "0000000000000000",
24899 => "0000000000000000",24900 => "0000000000000000",
24901 => "0000000000000000",24902 => "0000000000000000",
24903 => "0000000000000000",24904 => "0000000000000000",
24905 => "0000000000000000",24906 => "0000000000000000",
24907 => "0000000000000000",24908 => "0000000000000000",
24909 => "0000000000000000",24910 => "0000000000000000",
24911 => "0000000000000000",24912 => "0000000000000000",
24913 => "0000000000000000",24914 => "0000000000000000",
24915 => "0000000000000000",24916 => "0000000000000000",
24917 => "0000000000000000",24918 => "0000000000000000",
24919 => "0000000000000000",24920 => "0000000000000000",
24921 => "0000000000000000",24922 => "0000000000000000",
24923 => "0000000000000000",24924 => "0000000000000000",
24925 => "0000000000000000",24926 => "0000000000000000",
24927 => "0000000000000000",24928 => "0000000000000000",
24929 => "0000000000000000",24930 => "0000000000000000",
24931 => "0000000000000000",24932 => "0000000000000000",
24933 => "0000000000000000",24934 => "0000000000000000",
24935 => "0000000000000000",24936 => "0000000000000000",
24937 => "0000000000000000",24938 => "0000000000000000",
24939 => "0000000000000000",24940 => "0000000000000000",
24941 => "0000000000000000",24942 => "0000000000000000",
24943 => "0000000000000000",24944 => "0000000000000000",
24945 => "0000000000000000",24946 => "0000000000000000",
24947 => "0000000000000000",24948 => "0000000000000000",
24949 => "0000000000000000",24950 => "0000000000000000",
24951 => "0000000000000000",24952 => "0000000000000000",
24953 => "0000000000000000",24954 => "0000000000000000",
24955 => "0000000000000000",24956 => "0000000000000000",
24957 => "0000000000000000",24958 => "0000000000000000",
24959 => "0000000000000000",24960 => "0000000000000000",
24961 => "0000000000000000",24962 => "0000000000000000",
24963 => "0000000000000000",24964 => "0000000000000000",
24965 => "0000000000000000",24966 => "0000000000000000",
24967 => "0000000000000000",24968 => "0000000000000000",
24969 => "0000000000000000",24970 => "0000000000000000",
24971 => "0000000000000000",24972 => "0000000000000000",
24973 => "0000000000000000",24974 => "0000000000000000",
24975 => "0000000000000000",24976 => "0000000000000000",
24977 => "0000000000000000",24978 => "0000000000000000",
24979 => "0000000000000000",24980 => "0000000000000000",
24981 => "0000000000000000",24982 => "0000000000000000",
24983 => "0000000000000000",24984 => "0000000000000000",
24985 => "0000000000000000",24986 => "0000000000000000",
24987 => "0000000000000000",24988 => "0000000000000000",
24989 => "0000000000000000",24990 => "0000000000000000",
24991 => "0000000000000000",24992 => "0000000000000000",
24993 => "0000000000000000",24994 => "0000000000000000",
24995 => "0000000000000000",24996 => "0000000000000000",
24997 => "0000000000000000",24998 => "0000000000000000",
24999 => "0000000000000000",25000 => "0000000000000000",
25001 => "0000000000000000",25002 => "0000000000000000",
25003 => "0000000000000000",25004 => "0000000000000000",
25005 => "0000000000000000",25006 => "0000000000000000",
25007 => "0000000000000000",25008 => "0000000000000000",
25009 => "0000000000000000",25010 => "0000000000000000",
25011 => "0000000000000000",25012 => "0000000000000000",
25013 => "0000000000000000",25014 => "0000000000000000",
25015 => "0000000000000000",25016 => "0000000000000000",
25017 => "0000000000000000",25018 => "0000000000000000",
25019 => "0000000000000000",25020 => "0000000000000000",
25021 => "0000000000000000",25022 => "0000000000000000",
25023 => "0000000000000000",25024 => "0000000000000000",
25025 => "0000000000000000",25026 => "0000000000000000",
25027 => "0000000000000000",25028 => "0000000000000000",
25029 => "0000000000000000",25030 => "0000000000000000",
25031 => "0000000000000000",25032 => "0000000000000000",
25033 => "0000000000000000",25034 => "0000000000000000",
25035 => "0000000000000000",25036 => "0000000000000000",
25037 => "0000000000000000",25038 => "0000000000000000",
25039 => "0000000000000000",25040 => "0000000000000000",
25041 => "0000000000000000",25042 => "0000000000000000",
25043 => "0000000000000000",25044 => "0000000000000000",
25045 => "0000000000000000",25046 => "0000000000000000",
25047 => "0000000000000000",25048 => "0000000000000000",
25049 => "0000000000000000",25050 => "0000000000000000",
25051 => "0000000000000000",25052 => "0000000000000000",
25053 => "0000000000000000",25054 => "0000000000000000",
25055 => "0000000000000000",25056 => "0000000000000000",
25057 => "0000000000000000",25058 => "0000000000000000",
25059 => "0000000000000000",25060 => "0000000000000000",
25061 => "0000000000000000",25062 => "0000000000000000",
25063 => "0000000000000000",25064 => "0000000000000000",
25065 => "0000000000000000",25066 => "0000000000000000",
25067 => "0000000000000000",25068 => "0000000000000000",
25069 => "0000000000000000",25070 => "0000000000000000",
25071 => "0000000000000000",25072 => "0000000000000000",
25073 => "0000000000000000",25074 => "0000000000000000",
25075 => "0000000000000000",25076 => "0000000000000000",
25077 => "0000000000000000",25078 => "0000000000000000",
25079 => "0000000000000000",25080 => "0000000000000000",
25081 => "0000000000000000",25082 => "0000000000000000",
25083 => "0000000000000000",25084 => "0000000000000000",
25085 => "0000000000000000",25086 => "0000000000000000",
25087 => "0000000000000000",25088 => "0000000000000000",
25089 => "0000000000000000",25090 => "0000000000000000",
25091 => "0000000000000000",25092 => "0000000000000000",
25093 => "0000000000000000",25094 => "0000000000000000",
25095 => "0000000000000000",25096 => "0000000000000000",
25097 => "0000000000000000",25098 => "0000000000000000",
25099 => "0000000000000000",25100 => "0000000000000000",
25101 => "0000000000000000",25102 => "0000000000000000",
25103 => "0000000000000000",25104 => "0000000000000000",
25105 => "0000000000000000",25106 => "0000000000000000",
25107 => "0000000000000000",25108 => "0000000000000000",
25109 => "0000000000000000",25110 => "0000000000000000",
25111 => "0000000000000000",25112 => "0000000000000000",
25113 => "0000000000000000",25114 => "0000000000000000",
25115 => "0000000000000000",25116 => "0000000000000000",
25117 => "0000000000000000",25118 => "0000000000000000",
25119 => "0000000000000000",25120 => "0000000000000000",
25121 => "0000000000000000",25122 => "0000000000000000",
25123 => "0000000000000000",25124 => "0000000000000000",
25125 => "0000000000000000",25126 => "0000000000000000",
25127 => "0000000000000000",25128 => "0000000000000000",
25129 => "0000000000000000",25130 => "0000000000000000",
25131 => "0000000000000000",25132 => "0000000000000000",
25133 => "0000000000000000",25134 => "0000000000000000",
25135 => "0000000000000000",25136 => "0000000000000000",
25137 => "0000000000000000",25138 => "0000000000000000",
25139 => "0000000000000000",25140 => "0000000000000000",
25141 => "0000000000000000",25142 => "0000000000000000",
25143 => "0000000000000000",25144 => "0000000000000000",
25145 => "0000000000000000",25146 => "0000000000000000",
25147 => "0000000000000000",25148 => "0000000000000000",
25149 => "0000000000000000",25150 => "0000000000000000",
25151 => "0000000000000000",25152 => "0000000000000000",
25153 => "0000000000000000",25154 => "0000000000000000",
25155 => "0000000000000000",25156 => "0000000000000000",
25157 => "0000000000000000",25158 => "0000000000000000",
25159 => "0000000000000000",25160 => "0000000000000000",
25161 => "0000000000000000",25162 => "0000000000000000",
25163 => "0000000000000000",25164 => "0000000000000000",
25165 => "0000000000000000",25166 => "0000000000000000",
25167 => "0000000000000000",25168 => "0000000000000000",
25169 => "0000000000000000",25170 => "0000000000000000",
25171 => "0000000000000000",25172 => "0000000000000000",
25173 => "0000000000000000",25174 => "0000000000000000",
25175 => "0000000000000000",25176 => "0000000000000000",
25177 => "0000000000000000",25178 => "0000000000000000",
25179 => "0000000000000000",25180 => "0000000000000000",
25181 => "0000000000000000",25182 => "0000000000000000",
25183 => "0000000000000000",25184 => "0000000000000000",
25185 => "0000000000000000",25186 => "0000000000000000",
25187 => "0000000000000000",25188 => "0000000000000000",
25189 => "0000000000000000",25190 => "0000000000000000",
25191 => "0000000000000000",25192 => "0000000000000000",
25193 => "0000000000000000",25194 => "0000000000000000",
25195 => "0000000000000000",25196 => "0000000000000000",
25197 => "0000000000000000",25198 => "0000000000000000",
25199 => "0000000000000000",25200 => "0000000000000000",
25201 => "0000000000000000",25202 => "0000000000000000",
25203 => "0000000000000000",25204 => "0000000000000000",
25205 => "0000000000000000",25206 => "0000000000000000",
25207 => "0000000000000000",25208 => "0000000000000000",
25209 => "0000000000000000",25210 => "0000000000000000",
25211 => "0000000000000000",25212 => "0000000000000000",
25213 => "0000000000000000",25214 => "0000000000000000",
25215 => "0000000000000000",25216 => "0000000000000000",
25217 => "0000000000000000",25218 => "0000000000000000",
25219 => "0000000000000000",25220 => "0000000000000000",
25221 => "0000000000000000",25222 => "0000000000000000",
25223 => "0000000000000000",25224 => "0000000000000000",
25225 => "0000000000000000",25226 => "0000000000000000",
25227 => "0000000000000000",25228 => "0000000000000000",
25229 => "0000000000000000",25230 => "0000000000000000",
25231 => "0000000000000000",25232 => "0000000000000000",
25233 => "0000000000000000",25234 => "0000000000000000",
25235 => "0000000000000000",25236 => "0000000000000000",
25237 => "0000000000000000",25238 => "0000000000000000",
25239 => "0000000000000000",25240 => "0000000000000000",
25241 => "0000000000000000",25242 => "0000000000000000",
25243 => "0000000000000000",25244 => "0000000000000000",
25245 => "0000000000000000",25246 => "0000000000000000",
25247 => "0000000000000000",25248 => "0000000000000000",
25249 => "0000000000000000",25250 => "0000000000000000",
25251 => "0000000000000000",25252 => "0000000000000000",
25253 => "0000000000000000",25254 => "0000000000000000",
25255 => "0000000000000000",25256 => "0000000000000000",
25257 => "0000000000000000",25258 => "0000000000000000",
25259 => "0000000000000000",25260 => "0000000000000000",
25261 => "0000000000000000",25262 => "0000000000000000",
25263 => "0000000000000000",25264 => "0000000000000000",
25265 => "0000000000000000",25266 => "0000000000000000",
25267 => "0000000000000000",25268 => "0000000000000000",
25269 => "0000000000000000",25270 => "0000000000000000",
25271 => "0000000000000000",25272 => "0000000000000000",
25273 => "0000000000000000",25274 => "0000000000000000",
25275 => "0000000000000000",25276 => "0000000000000000",
25277 => "0000000000000000",25278 => "0000000000000000",
25279 => "0000000000000000",25280 => "0000000000000000",
25281 => "0000000000000000",25282 => "0000000000000000",
25283 => "0000000000000000",25284 => "0000000000000000",
25285 => "0000000000000000",25286 => "0000000000000000",
25287 => "0000000000000000",25288 => "0000000000000000",
25289 => "0000000000000000",25290 => "0000000000000000",
25291 => "0000000000000000",25292 => "0000000000000000",
25293 => "0000000000000000",25294 => "0000000000000000",
25295 => "0000000000000000",25296 => "0000000000000000",
25297 => "0000000000000000",25298 => "0000000000000000",
25299 => "0000000000000000",25300 => "0000000000000000",
25301 => "0000000000000000",25302 => "0000000000000000",
25303 => "0000000000000000",25304 => "0000000000000000",
25305 => "0000000000000000",25306 => "0000000000000000",
25307 => "0000000000000000",25308 => "0000000000000000",
25309 => "0000000000000000",25310 => "0000000000000000",
25311 => "0000000000000000",25312 => "0000000000000000",
25313 => "0000000000000000",25314 => "0000000000000000",
25315 => "0000000000000000",25316 => "0000000000000000",
25317 => "0000000000000000",25318 => "0000000000000000",
25319 => "0000000000000000",25320 => "0000000000000000",
25321 => "0000000000000000",25322 => "0000000000000000",
25323 => "0000000000000000",25324 => "0000000000000000",
25325 => "0000000000000000",25326 => "0000000000000000",
25327 => "0000000000000000",25328 => "0000000000000000",
25329 => "0000000000000000",25330 => "0000000000000000",
25331 => "0000000000000000",25332 => "0000000000000000",
25333 => "0000000000000000",25334 => "0000000000000000",
25335 => "0000000000000000",25336 => "0000000000000000",
25337 => "0000000000000000",25338 => "0000000000000000",
25339 => "0000000000000000",25340 => "0000000000000000",
25341 => "0000000000000000",25342 => "0000000000000000",
25343 => "0000000000000000",25344 => "0000000000000000",
25345 => "0000000000000000",25346 => "0000000000000000",
25347 => "0000000000000000",25348 => "0000000000000000",
25349 => "0000000000000000",25350 => "0000000000000000",
25351 => "0000000000000000",25352 => "0000000000000000",
25353 => "0000000000000000",25354 => "0000000000000000",
25355 => "0000000000000000",25356 => "0000000000000000",
25357 => "0000000000000000",25358 => "0000000000000000",
25359 => "0000000000000000",25360 => "0000000000000000",
25361 => "0000000000000000",25362 => "0000000000000000",
25363 => "0000000000000000",25364 => "0000000000000000",
25365 => "0000000000000000",25366 => "0000000000000000",
25367 => "0000000000000000",25368 => "0000000000000000",
25369 => "0000000000000000",25370 => "0000000000000000",
25371 => "0000000000000000",25372 => "0000000000000000",
25373 => "0000000000000000",25374 => "0000000000000000",
25375 => "0000000000000000",25376 => "0000000000000000",
25377 => "0000000000000000",25378 => "0000000000000000",
25379 => "0000000000000000",25380 => "0000000000000000",
25381 => "0000000000000000",25382 => "0000000000000000",
25383 => "0000000000000000",25384 => "0000000000000000",
25385 => "0000000000000000",25386 => "0000000000000000",
25387 => "0000000000000000",25388 => "0000000000000000",
25389 => "0000000000000000",25390 => "0000000000000000",
25391 => "0000000000000000",25392 => "0000000000000000",
25393 => "0000000000000000",25394 => "0000000000000000",
25395 => "0000000000000000",25396 => "0000000000000000",
25397 => "0000000000000000",25398 => "0000000000000000",
25399 => "0000000000000000",25400 => "0000000000000000",
25401 => "0000000000000000",25402 => "0000000000000000",
25403 => "0000000000000000",25404 => "0000000000000000",
25405 => "0000000000000000",25406 => "0000000000000000",
25407 => "0000000000000000",25408 => "0000000000000000",
25409 => "0000000000000000",25410 => "0000000000000000",
25411 => "0000000000000000",25412 => "0000000000000000",
25413 => "0000000000000000",25414 => "0000000000000000",
25415 => "0000000000000000",25416 => "0000000000000000",
25417 => "0000000000000000",25418 => "0000000000000000",
25419 => "0000000000000000",25420 => "0000000000000000",
25421 => "0000000000000000",25422 => "0000000000000000",
25423 => "0000000000000000",25424 => "0000000000000000",
25425 => "0000000000000000",25426 => "0000000000000000",
25427 => "0000000000000000",25428 => "0000000000000000",
25429 => "0000000000000000",25430 => "0000000000000000",
25431 => "0000000000000000",25432 => "0000000000000000",
25433 => "0000000000000000",25434 => "0000000000000000",
25435 => "0000000000000000",25436 => "0000000000000000",
25437 => "0000000000000000",25438 => "0000000000000000",
25439 => "0000000000000000",25440 => "0000000000000000",
25441 => "0000000000000000",25442 => "0000000000000000",
25443 => "0000000000000000",25444 => "0000000000000000",
25445 => "0000000000000000",25446 => "0000000000000000",
25447 => "0000000000000000",25448 => "0000000000000000",
25449 => "0000000000000000",25450 => "0000000000000000",
25451 => "0000000000000000",25452 => "0000000000000000",
25453 => "0000000000000000",25454 => "0000000000000000",
25455 => "0000000000000000",25456 => "0000000000000000",
25457 => "0000000000000000",25458 => "0000000000000000",
25459 => "0000000000000000",25460 => "0000000000000000",
25461 => "0000000000000000",25462 => "0000000000000000",
25463 => "0000000000000000",25464 => "0000000000000000",
25465 => "0000000000000000",25466 => "0000000000000000",
25467 => "0000000000000000",25468 => "0000000000000000",
25469 => "0000000000000000",25470 => "0000000000000000",
25471 => "0000000000000000",25472 => "0000000000000000",
25473 => "0000000000000000",25474 => "0000000000000000",
25475 => "0000000000000000",25476 => "0000000000000000",
25477 => "0000000000000000",25478 => "0000000000000000",
25479 => "0000000000000000",25480 => "0000000000000000",
25481 => "0000000000000000",25482 => "0000000000000000",
25483 => "0000000000000000",25484 => "0000000000000000",
25485 => "0000000000000000",25486 => "0000000000000000",
25487 => "0000000000000000",25488 => "0000000000000000",
25489 => "0000000000000000",25490 => "0000000000000000",
25491 => "0000000000000000",25492 => "0000000000000000",
25493 => "0000000000000000",25494 => "0000000000000000",
25495 => "0000000000000000",25496 => "0000000000000000",
25497 => "0000000000000000",25498 => "0000000000000000",
25499 => "0000000000000000",25500 => "0000000000000000",
25501 => "0000000000000000",25502 => "0000000000000000",
25503 => "0000000000000000",25504 => "0000000000000000",
25505 => "0000000000000000",25506 => "0000000000000000",
25507 => "0000000000000000",25508 => "0000000000000000",
25509 => "0000000000000000",25510 => "0000000000000000",
25511 => "0000000000000000",25512 => "0000000000000000",
25513 => "0000000000000000",25514 => "0000000000000000",
25515 => "0000000000000000",25516 => "0000000000000000",
25517 => "0000000000000000",25518 => "0000000000000000",
25519 => "0000000000000000",25520 => "0000000000000000",
25521 => "0000000000000000",25522 => "0000000000000000",
25523 => "0000000000000000",25524 => "0000000000000000",
25525 => "0000000000000000",25526 => "0000000000000000",
25527 => "0000000000000000",25528 => "0000000000000000",
25529 => "0000000000000000",25530 => "0000000000000000",
25531 => "0000000000000000",25532 => "0000000000000000",
25533 => "0000000000000000",25534 => "0000000000000000",
25535 => "0000000000000000",25536 => "0000000000000000",
25537 => "0000000000000000",25538 => "0000000000000000",
25539 => "0000000000000000",25540 => "0000000000000000",
25541 => "0000000000000000",25542 => "0000000000000000",
25543 => "0000000000000000",25544 => "0000000000000000",
25545 => "0000000000000000",25546 => "0000000000000000",
25547 => "0000000000000000",25548 => "0000000000000000",
25549 => "0000000000000000",25550 => "0000000000000000",
25551 => "0000000000000000",25552 => "0000000000000000",
25553 => "0000000000000000",25554 => "0000000000000000",
25555 => "0000000000000000",25556 => "0000000000000000",
25557 => "0000000000000000",25558 => "0000000000000000",
25559 => "0000000000000000",25560 => "0000000000000000",
25561 => "0000000000000000",25562 => "0000000000000000",
25563 => "0000000000000000",25564 => "0000000000000000",
25565 => "0000000000000000",25566 => "0000000000000000",
25567 => "0000000000000000",25568 => "0000000000000000",
25569 => "0000000000000000",25570 => "0000000000000000",
25571 => "0000000000000000",25572 => "0000000000000000",
25573 => "0000000000000000",25574 => "0000000000000000",
25575 => "0000000000000000",25576 => "0000000000000000",
25577 => "0000000000000000",25578 => "0000000000000000",
25579 => "0000000000000000",25580 => "0000000000000000",
25581 => "0000000000000000",25582 => "0000000000000000",
25583 => "0000000000000000",25584 => "0000000000000000",
25585 => "0000000000000000",25586 => "0000000000000000",
25587 => "0000000000000000",25588 => "0000000000000000",
25589 => "0000000000000000",25590 => "0000000000000000",
25591 => "0000000000000000",25592 => "0000000000000000",
25593 => "0000000000000000",25594 => "0000000000000000",
25595 => "0000000000000000",25596 => "0000000000000000",
25597 => "0000000000000000",25598 => "0000000000000000",
25599 => "0000000000000000",25600 => "0000000000000000",
25601 => "0000000000000000",25602 => "0000000000000000",
25603 => "0000000000000000",25604 => "0000000000000000",
25605 => "0000000000000000",25606 => "0000000000000000",
25607 => "0000000000000000",25608 => "0000000000000000",
25609 => "0000000000000000",25610 => "0000000000000000",
25611 => "0000000000000000",25612 => "0000000000000000",
25613 => "0000000000000000",25614 => "0000000000000000",
25615 => "0000000000000000",25616 => "0000000000000000",
25617 => "0000000000000000",25618 => "0000000000000000",
25619 => "0000000000000000",25620 => "0000000000000000",
25621 => "0000000000000000",25622 => "0000000000000000",
25623 => "0000000000000000",25624 => "0000000000000000",
25625 => "0000000000000000",25626 => "0000000000000000",
25627 => "0000000000000000",25628 => "0000000000000000",
25629 => "0000000000000000",25630 => "0000000000000000",
25631 => "0000000000000000",25632 => "0000000000000000",
25633 => "0000000000000000",25634 => "0000000000000000",
25635 => "0000000000000000",25636 => "0000000000000000",
25637 => "0000000000000000",25638 => "0000000000000000",
25639 => "0000000000000000",25640 => "0000000000000000",
25641 => "0000000000000000",25642 => "0000000000000000",
25643 => "0000000000000000",25644 => "0000000000000000",
25645 => "0000000000000000",25646 => "0000000000000000",
25647 => "0000000000000000",25648 => "0000000000000000",
25649 => "0000000000000000",25650 => "0000000000000000",
25651 => "0000000000000000",25652 => "0000000000000000",
25653 => "0000000000000000",25654 => "0000000000000000",
25655 => "0000000000000000",25656 => "0000000000000000",
25657 => "0000000000000000",25658 => "0000000000000000",
25659 => "0000000000000000",25660 => "0000000000000000",
25661 => "0000000000000000",25662 => "0000000000000000",
25663 => "0000000000000000",25664 => "0000000000000000",
25665 => "0000000000000000",25666 => "0000000000000000",
25667 => "0000000000000000",25668 => "0000000000000000",
25669 => "0000000000000000",25670 => "0000000000000000",
25671 => "0000000000000000",25672 => "0000000000000000",
25673 => "0000000000000000",25674 => "0000000000000000",
25675 => "0000000000000000",25676 => "0000000000000000",
25677 => "0000000000000000",25678 => "0000000000000000",
25679 => "0000000000000000",25680 => "0000000000000000",
25681 => "0000000000000000",25682 => "0000000000000000",
25683 => "0000000000000000",25684 => "0000000000000000",
25685 => "0000000000000000",25686 => "0000000000000000",
25687 => "0000000000000000",25688 => "0000000000000000",
25689 => "0000000000000000",25690 => "0000000000000000",
25691 => "0000000000000000",25692 => "0000000000000000",
25693 => "0000000000000000",25694 => "0000000000000000",
25695 => "0000000000000000",25696 => "0000000000000000",
25697 => "0000000000000000",25698 => "0000000000000000",
25699 => "0000000000000000",25700 => "0000000000000000",
25701 => "0000000000000000",25702 => "0000000000000000",
25703 => "0000000000000000",25704 => "0000000000000000",
25705 => "0000000000000000",25706 => "0000000000000000",
25707 => "0000000000000000",25708 => "0000000000000000",
25709 => "0000000000000000",25710 => "0000000000000000",
25711 => "0000000000000000",25712 => "0000000000000000",
25713 => "0000000000000000",25714 => "0000000000000000",
25715 => "0000000000000000",25716 => "0000000000000000",
25717 => "0000000000000000",25718 => "0000000000000000",
25719 => "0000000000000000",25720 => "0000000000000000",
25721 => "0000000000000000",25722 => "0000000000000000",
25723 => "0000000000000000",25724 => "0000000000000000",
25725 => "0000000000000000",25726 => "0000000000000000",
25727 => "0000000000000000",25728 => "0000000000000000",
25729 => "0000000000000000",25730 => "0000000000000000",
25731 => "0000000000000000",25732 => "0000000000000000",
25733 => "0000000000000000",25734 => "0000000000000000",
25735 => "0000000000000000",25736 => "0000000000000000",
25737 => "0000000000000000",25738 => "0000000000000000",
25739 => "0000000000000000",25740 => "0000000000000000",
25741 => "0000000000000000",25742 => "0000000000000000",
25743 => "0000000000000000",25744 => "0000000000000000",
25745 => "0000000000000000",25746 => "0000000000000000",
25747 => "0000000000000000",25748 => "0000000000000000",
25749 => "0000000000000000",25750 => "0000000000000000",
25751 => "0000000000000000",25752 => "0000000000000000",
25753 => "0000000000000000",25754 => "0000000000000000",
25755 => "0000000000000000",25756 => "0000000000000000",
25757 => "0000000000000000",25758 => "0000000000000000",
25759 => "0000000000000000",25760 => "0000000000000000",
25761 => "0000000000000000",25762 => "0000000000000000",
25763 => "0000000000000000",25764 => "0000000000000000",
25765 => "0000000000000000",25766 => "0000000000000000",
25767 => "0000000000000000",25768 => "0000000000000000",
25769 => "0000000000000000",25770 => "0000000000000000",
25771 => "0000000000000000",25772 => "0000000000000000",
25773 => "0000000000000000",25774 => "0000000000000000",
25775 => "0000000000000000",25776 => "0000000000000000",
25777 => "0000000000000000",25778 => "0000000000000000",
25779 => "0000000000000000",25780 => "0000000000000000",
25781 => "0000000000000000",25782 => "0000000000000000",
25783 => "0000000000000000",25784 => "0000000000000000",
25785 => "0000000000000000",25786 => "0000000000000000",
25787 => "0000000000000000",25788 => "0000000000000000",
25789 => "0000000000000000",25790 => "0000000000000000",
25791 => "0000000000000000",25792 => "0000000000000000",
25793 => "0000000000000000",25794 => "0000000000000000",
25795 => "0000000000000000",25796 => "0000000000000000",
25797 => "0000000000000000",25798 => "0000000000000000",
25799 => "0000000000000000",25800 => "0000000000000000",
25801 => "0000000000000000",25802 => "0000000000000000",
25803 => "0000000000000000",25804 => "0000000000000000",
25805 => "0000000000000000",25806 => "0000000000000000",
25807 => "0000000000000000",25808 => "0000000000000000",
25809 => "0000000000000000",25810 => "0000000000000000",
25811 => "0000000000000000",25812 => "0000000000000000",
25813 => "0000000000000000",25814 => "0000000000000000",
25815 => "0000000000000000",25816 => "0000000000000000",
25817 => "0000000000000000",25818 => "0000000000000000",
25819 => "0000000000000000",25820 => "0000000000000000",
25821 => "0000000000000000",25822 => "0000000000000000",
25823 => "0000000000000000",25824 => "0000000000000000",
25825 => "0000000000000000",25826 => "0000000000000000",
25827 => "0000000000000000",25828 => "0000000000000000",
25829 => "0000000000000000",25830 => "0000000000000000",
25831 => "0000000000000000",25832 => "0000000000000000",
25833 => "0000000000000000",25834 => "0000000000000000",
25835 => "0000000000000000",25836 => "0000000000000000",
25837 => "0000000000000000",25838 => "0000000000000000",
25839 => "0000000000000000",25840 => "0000000000000000",
25841 => "0000000000000000",25842 => "0000000000000000",
25843 => "0000000000000000",25844 => "0000000000000000",
25845 => "0000000000000000",25846 => "0000000000000000",
25847 => "0000000000000000",25848 => "0000000000000000",
25849 => "0000000000000000",25850 => "0000000000000000",
25851 => "0000000000000000",25852 => "0000000000000000",
25853 => "0000000000000000",25854 => "0000000000000000",
25855 => "0000000000000000",25856 => "0000000000000000",
25857 => "0000000000000000",25858 => "0000000000000000",
25859 => "0000000000000000",25860 => "0000000000000000",
25861 => "0000000000000000",25862 => "0000000000000000",
25863 => "0000000000000000",25864 => "0000000000000000",
25865 => "0000000000000000",25866 => "0000000000000000",
25867 => "0000000000000000",25868 => "0000000000000000",
25869 => "0000000000000000",25870 => "0000000000000000",
25871 => "0000000000000000",25872 => "0000000000000000",
25873 => "0000000000000000",25874 => "0000000000000000",
25875 => "0000000000000000",25876 => "0000000000000000",
25877 => "0000000000000000",25878 => "0000000000000000",
25879 => "0000000000000000",25880 => "0000000000000000",
25881 => "0000000000000000",25882 => "0000000000000000",
25883 => "0000000000000000",25884 => "0000000000000000",
25885 => "0000000000000000",25886 => "0000000000000000",
25887 => "0000000000000000",25888 => "0000000000000000",
25889 => "0000000000000000",25890 => "0000000000000000",
25891 => "0000000000000000",25892 => "0000000000000000",
25893 => "0000000000000000",25894 => "0000000000000000",
25895 => "0000000000000000",25896 => "0000000000000000",
25897 => "0000000000000000",25898 => "0000000000000000",
25899 => "0000000000000000",25900 => "0000000000000000",
25901 => "0000000000000000",25902 => "0000000000000000",
25903 => "0000000000000000",25904 => "0000000000000000",
25905 => "0000000000000000",25906 => "0000000000000000",
25907 => "0000000000000000",25908 => "0000000000000000",
25909 => "0000000000000000",25910 => "0000000000000000",
25911 => "0000000000000000",25912 => "0000000000000000",
25913 => "0000000000000000",25914 => "0000000000000000",
25915 => "0000000000000000",25916 => "0000000000000000",
25917 => "0000000000000000",25918 => "0000000000000000",
25919 => "0000000000000000",25920 => "0000000000000000",
25921 => "0000000000000000",25922 => "0000000000000000",
25923 => "0000000000000000",25924 => "0000000000000000",
25925 => "0000000000000000",25926 => "0000000000000000",
25927 => "0000000000000000",25928 => "0000000000000000",
25929 => "0000000000000000",25930 => "0000000000000000",
25931 => "0000000000000000",25932 => "0000000000000000",
25933 => "0000000000000000",25934 => "0000000000000000",
25935 => "0000000000000000",25936 => "0000000000000000",
25937 => "0000000000000000",25938 => "0000000000000000",
25939 => "0000000000000000",25940 => "0000000000000000",
25941 => "0000000000000000",25942 => "0000000000000000",
25943 => "0000000000000000",25944 => "0000000000000000",
25945 => "0000000000000000",25946 => "0000000000000000",
25947 => "0000000000000000",25948 => "0000000000000000",
25949 => "0000000000000000",25950 => "0000000000000000",
25951 => "0000000000000000",25952 => "0000000000000000",
25953 => "0000000000000000",25954 => "0000000000000000",
25955 => "0000000000000000",25956 => "0000000000000000",
25957 => "0000000000000000",25958 => "0000000000000000",
25959 => "0000000000000000",25960 => "0000000000000000",
25961 => "0000000000000000",25962 => "0000000000000000",
25963 => "0000000000000000",25964 => "0000000000000000",
25965 => "0000000000000000",25966 => "0000000000000000",
25967 => "0000000000000000",25968 => "0000000000000000",
25969 => "0000000000000000",25970 => "0000000000000000",
25971 => "0000000000000000",25972 => "0000000000000000",
25973 => "0000000000000000",25974 => "0000000000000000",
25975 => "0000000000000000",25976 => "0000000000000000",
25977 => "0000000000000000",25978 => "0000000000000000",
25979 => "0000000000000000",25980 => "0000000000000000",
25981 => "0000000000000000",25982 => "0000000000000000",
25983 => "0000000000000000",25984 => "0000000000000000",
25985 => "0000000000000000",25986 => "0000000000000000",
25987 => "0000000000000000",25988 => "0000000000000000",
25989 => "0000000000000000",25990 => "0000000000000000",
25991 => "0000000000000000",25992 => "0000000000000000",
25993 => "0000000000000000",25994 => "0000000000000000",
25995 => "0000000000000000",25996 => "0000000000000000",
25997 => "0000000000000000",25998 => "0000000000000000",
25999 => "0000000000000000",26000 => "0000000000000000",
26001 => "0000000000000000",26002 => "0000000000000000",
26003 => "0000000000000000",26004 => "0000000000000000",
26005 => "0000000000000000",26006 => "0000000000000000",
26007 => "0000000000000000",26008 => "0000000000000000",
26009 => "0000000000000000",26010 => "0000000000000000",
26011 => "0000000000000000",26012 => "0000000000000000",
26013 => "0000000000000000",26014 => "0000000000000000",
26015 => "0000000000000000",26016 => "0000000000000000",
26017 => "0000000000000000",26018 => "0000000000000000",
26019 => "0000000000000000",26020 => "0000000000000000",
26021 => "0000000000000000",26022 => "0000000000000000",
26023 => "0000000000000000",26024 => "0000000000000000",
26025 => "0000000000000000",26026 => "0000000000000000",
26027 => "0000000000000000",26028 => "0000000000000000",
26029 => "0000000000000000",26030 => "0000000000000000",
26031 => "0000000000000000",26032 => "0000000000000000",
26033 => "0000000000000000",26034 => "0000000000000000",
26035 => "0000000000000000",26036 => "0000000000000000",
26037 => "0000000000000000",26038 => "0000000000000000",
26039 => "0000000000000000",26040 => "0000000000000000",
26041 => "0000000000000000",26042 => "0000000000000000",
26043 => "0000000000000000",26044 => "0000000000000000",
26045 => "0000000000000000",26046 => "0000000000000000",
26047 => "0000000000000000",26048 => "0000000000000000",
26049 => "0000000000000000",26050 => "0000000000000000",
26051 => "0000000000000000",26052 => "0000000000000000",
26053 => "0000000000000000",26054 => "0000000000000000",
26055 => "0000000000000000",26056 => "0000000000000000",
26057 => "0000000000000000",26058 => "0000000000000000",
26059 => "0000000000000000",26060 => "0000000000000000",
26061 => "0000000000000000",26062 => "0000000000000000",
26063 => "0000000000000000",26064 => "0000000000000000",
26065 => "0000000000000000",26066 => "0000000000000000",
26067 => "0000000000000000",26068 => "0000000000000000",
26069 => "0000000000000000",26070 => "0000000000000000",
26071 => "0000000000000000",26072 => "0000000000000000",
26073 => "0000000000000000",26074 => "0000000000000000",
26075 => "0000000000000000",26076 => "0000000000000000",
26077 => "0000000000000000",26078 => "0000000000000000",
26079 => "0000000000000000",26080 => "0000000000000000",
26081 => "0000000000000000",26082 => "0000000000000000",
26083 => "0000000000000000",26084 => "0000000000000000",
26085 => "0000000000000000",26086 => "0000000000000000",
26087 => "0000000000000000",26088 => "0000000000000000",
26089 => "0000000000000000",26090 => "0000000000000000",
26091 => "0000000000000000",26092 => "0000000000000000",
26093 => "0000000000000000",26094 => "0000000000000000",
26095 => "0000000000000000",26096 => "0000000000000000",
26097 => "0000000000000000",26098 => "0000000000000000",
26099 => "0000000000000000",26100 => "0000000000000000",
26101 => "0000000000000000",26102 => "0000000000000000",
26103 => "0000000000000000",26104 => "0000000000000000",
26105 => "0000000000000000",26106 => "0000000000000000",
26107 => "0000000000000000",26108 => "0000000000000000",
26109 => "0000000000000000",26110 => "0000000000000000",
26111 => "0000000000000000",26112 => "0000000000000000",
26113 => "0000000000000000",26114 => "0000000000000000",
26115 => "0000000000000000",26116 => "0000000000000000",
26117 => "0000000000000000",26118 => "0000000000000000",
26119 => "0000000000000000",26120 => "0000000000000000",
26121 => "0000000000000000",26122 => "0000000000000000",
26123 => "0000000000000000",26124 => "0000000000000000",
26125 => "0000000000000000",26126 => "0000000000000000",
26127 => "0000000000000000",26128 => "0000000000000000",
26129 => "0000000000000000",26130 => "0000000000000000",
26131 => "0000000000000000",26132 => "0000000000000000",
26133 => "0000000000000000",26134 => "0000000000000000",
26135 => "0000000000000000",26136 => "0000000000000000",
26137 => "0000000000000000",26138 => "0000000000000000",
26139 => "0000000000000000",26140 => "0000000000000000",
26141 => "0000000000000000",26142 => "0000000000000000",
26143 => "0000000000000000",26144 => "0000000000000000",
26145 => "0000000000000000",26146 => "0000000000000000",
26147 => "0000000000000000",26148 => "0000000000000000",
26149 => "0000000000000000",26150 => "0000000000000000",
26151 => "0000000000000000",26152 => "0000000000000000",
26153 => "0000000000000000",26154 => "0000000000000000",
26155 => "0000000000000000",26156 => "0000000000000000",
26157 => "0000000000000000",26158 => "0000000000000000",
26159 => "0000000000000000",26160 => "0000000000000000",
26161 => "0000000000000000",26162 => "0000000000000000",
26163 => "0000000000000000",26164 => "0000000000000000",
26165 => "0000000000000000",26166 => "0000000000000000",
26167 => "0000000000000000",26168 => "0000000000000000",
26169 => "0000000000000000",26170 => "0000000000000000",
26171 => "0000000000000000",26172 => "0000000000000000",
26173 => "0000000000000000",26174 => "0000000000000000",
26175 => "0000000000000000",26176 => "0000000000000000",
26177 => "0000000000000000",26178 => "0000000000000000",
26179 => "0000000000000000",26180 => "0000000000000000",
26181 => "0000000000000000",26182 => "0000000000000000",
26183 => "0000000000000000",26184 => "0000000000000000",
26185 => "0000000000000000",26186 => "0000000000000000",
26187 => "0000000000000000",26188 => "0000000000000000",
26189 => "0000000000000000",26190 => "0000000000000000",
26191 => "0000000000000000",26192 => "0000000000000000",
26193 => "0000000000000000",26194 => "0000000000000000",
26195 => "0000000000000000",26196 => "0000000000000000",
26197 => "0000000000000000",26198 => "0000000000000000",
26199 => "0000000000000000",26200 => "0000000000000000",
26201 => "0000000000000000",26202 => "0000000000000000",
26203 => "0000000000000000",26204 => "0000000000000000",
26205 => "0000000000000000",26206 => "0000000000000000",
26207 => "0000000000000000",26208 => "0000000000000000",
26209 => "0000000000000000",26210 => "0000000000000000",
26211 => "0000000000000000",26212 => "0000000000000000",
26213 => "0000000000000000",26214 => "0000000000000000",
26215 => "0000000000000000",26216 => "0000000000000000",
26217 => "0000000000000000",26218 => "0000000000000000",
26219 => "0000000000000000",26220 => "0000000000000000",
26221 => "0000000000000000",26222 => "0000000000000000",
26223 => "0000000000000000",26224 => "0000000000000000",
26225 => "0000000000000000",26226 => "0000000000000000",
26227 => "0000000000000000",26228 => "0000000000000000",
26229 => "0000000000000000",26230 => "0000000000000000",
26231 => "0000000000000000",26232 => "0000000000000000",
26233 => "0000000000000000",26234 => "0000000000000000",
26235 => "0000000000000000",26236 => "0000000000000000",
26237 => "0000000000000000",26238 => "0000000000000000",
26239 => "0000000000000000",26240 => "0000000000000000",
26241 => "0000000000000000",26242 => "0000000000000000",
26243 => "0000000000000000",26244 => "0000000000000000",
26245 => "0000000000000000",26246 => "0000000000000000",
26247 => "0000000000000000",26248 => "0000000000000000",
26249 => "0000000000000000",26250 => "0000000000000000",
26251 => "0000000000000000",26252 => "0000000000000000",
26253 => "0000000000000000",26254 => "0000000000000000",
26255 => "0000000000000000",26256 => "0000000000000000",
26257 => "0000000000000000",26258 => "0000000000000000",
26259 => "0000000000000000",26260 => "0000000000000000",
26261 => "0000000000000000",26262 => "0000000000000000",
26263 => "0000000000000000",26264 => "0000000000000000",
26265 => "0000000000000000",26266 => "0000000000000000",
26267 => "0000000000000000",26268 => "0000000000000000",
26269 => "0000000000000000",26270 => "0000000000000000",
26271 => "0000000000000000",26272 => "0000000000000000",
26273 => "0000000000000000",26274 => "0000000000000000",
26275 => "0000000000000000",26276 => "0000000000000000",
26277 => "0000000000000000",26278 => "0000000000000000",
26279 => "0000000000000000",26280 => "0000000000000000",
26281 => "0000000000000000",26282 => "0000000000000000",
26283 => "0000000000000000",26284 => "0000000000000000",
26285 => "0000000000000000",26286 => "0000000000000000",
26287 => "0000000000000000",26288 => "0000000000000000",
26289 => "0000000000000000",26290 => "0000000000000000",
26291 => "0000000000000000",26292 => "0000000000000000",
26293 => "0000000000000000",26294 => "0000000000000000",
26295 => "0000000000000000",26296 => "0000000000000000",
26297 => "0000000000000000",26298 => "0000000000000000",
26299 => "0000000000000000",26300 => "0000000000000000",
26301 => "0000000000000000",26302 => "0000000000000000",
26303 => "0000000000000000",26304 => "0000000000000000",
26305 => "0000000000000000",26306 => "0000000000000000",
26307 => "0000000000000000",26308 => "0000000000000000",
26309 => "0000000000000000",26310 => "0000000000000000",
26311 => "0000000000000000",26312 => "0000000000000000",
26313 => "0000000000000000",26314 => "0000000000000000",
26315 => "0000000000000000",26316 => "0000000000000000",
26317 => "0000000000000000",26318 => "0000000000000000",
26319 => "0000000000000000",26320 => "0000000000000000",
26321 => "0000000000000000",26322 => "0000000000000000",
26323 => "0000000000000000",26324 => "0000000000000000",
26325 => "0000000000000000",26326 => "0000000000000000",
26327 => "0000000000000000",26328 => "0000000000000000",
26329 => "0000000000000000",26330 => "0000000000000000",
26331 => "0000000000000000",26332 => "0000000000000000",
26333 => "0000000000000000",26334 => "0000000000000000",
26335 => "0000000000000000",26336 => "0000000000000000",
26337 => "0000000000000000",26338 => "0000000000000000",
26339 => "0000000000000000",26340 => "0000000000000000",
26341 => "0000000000000000",26342 => "0000000000000000",
26343 => "0000000000000000",26344 => "0000000000000000",
26345 => "0000000000000000",26346 => "0000000000000000",
26347 => "0000000000000000",26348 => "0000000000000000",
26349 => "0000000000000000",26350 => "0000000000000000",
26351 => "0000000000000000",26352 => "0000000000000000",
26353 => "0000000000000000",26354 => "0000000000000000",
26355 => "0000000000000000",26356 => "0000000000000000",
26357 => "0000000000000000",26358 => "0000000000000000",
26359 => "0000000000000000",26360 => "0000000000000000",
26361 => "0000000000000000",26362 => "0000000000000000",
26363 => "0000000000000000",26364 => "0000000000000000",
26365 => "0000000000000000",26366 => "0000000000000000",
26367 => "0000000000000000",26368 => "0000000000000000",
26369 => "0000000000000000",26370 => "0000000000000000",
26371 => "0000000000000000",26372 => "0000000000000000",
26373 => "0000000000000000",26374 => "0000000000000000",
26375 => "0000000000000000",26376 => "0000000000000000",
26377 => "0000000000000000",26378 => "0000000000000000",
26379 => "0000000000000000",26380 => "0000000000000000",
26381 => "0000000000000000",26382 => "0000000000000000",
26383 => "0000000000000000",26384 => "0000000000000000",
26385 => "0000000000000000",26386 => "0000000000000000",
26387 => "0000000000000000",26388 => "0000000000000000",
26389 => "0000000000000000",26390 => "0000000000000000",
26391 => "0000000000000000",26392 => "0000000000000000",
26393 => "0000000000000000",26394 => "0000000000000000",
26395 => "0000000000000000",26396 => "0000000000000000",
26397 => "0000000000000000",26398 => "0000000000000000",
26399 => "0000000000000000",26400 => "0000000000000000",
26401 => "0000000000000000",26402 => "0000000000000000",
26403 => "0000000000000000",26404 => "0000000000000000",
26405 => "0000000000000000",26406 => "0000000000000000",
26407 => "0000000000000000",26408 => "0000000000000000",
26409 => "0000000000000000",26410 => "0000000000000000",
26411 => "0000000000000000",26412 => "0000000000000000",
26413 => "0000000000000000",26414 => "0000000000000000",
26415 => "0000000000000000",26416 => "0000000000000000",
26417 => "0000000000000000",26418 => "0000000000000000",
26419 => "0000000000000000",26420 => "0000000000000000",
26421 => "0000000000000000",26422 => "0000000000000000",
26423 => "0000000000000000",26424 => "0000000000000000",
26425 => "0000000000000000",26426 => "0000000000000000",
26427 => "0000000000000000",26428 => "0000000000000000",
26429 => "0000000000000000",26430 => "0000000000000000",
26431 => "0000000000000000",26432 => "0000000000000000",
26433 => "0000000000000000",26434 => "0000000000000000",
26435 => "0000000000000000",26436 => "0000000000000000",
26437 => "0000000000000000",26438 => "0000000000000000",
26439 => "0000000000000000",26440 => "0000000000000000",
26441 => "0000000000000000",26442 => "0000000000000000",
26443 => "0000000000000000",26444 => "0000000000000000",
26445 => "0000000000000000",26446 => "0000000000000000",
26447 => "0000000000000000",26448 => "0000000000000000",
26449 => "0000000000000000",26450 => "0000000000000000",
26451 => "0000000000000000",26452 => "0000000000000000",
26453 => "0000000000000000",26454 => "0000000000000000",
26455 => "0000000000000000",26456 => "0000000000000000",
26457 => "0000000000000000",26458 => "0000000000000000",
26459 => "0000000000000000",26460 => "0000000000000000",
26461 => "0000000000000000",26462 => "0000000000000000",
26463 => "0000000000000000",26464 => "0000000000000000",
26465 => "0000000000000000",26466 => "0000000000000000",
26467 => "0000000000000000",26468 => "0000000000000000",
26469 => "0000000000000000",26470 => "0000000000000000",
26471 => "0000000000000000",26472 => "0000000000000000",
26473 => "0000000000000000",26474 => "0000000000000000",
26475 => "0000000000000000",26476 => "0000000000000000",
26477 => "0000000000000000",26478 => "0000000000000000",
26479 => "0000000000000000",26480 => "0000000000000000",
26481 => "0000000000000000",26482 => "0000000000000000",
26483 => "0000000000000000",26484 => "0000000000000000",
26485 => "0000000000000000",26486 => "0000000000000000",
26487 => "0000000000000000",26488 => "0000000000000000",
26489 => "0000000000000000",26490 => "0000000000000000",
26491 => "0000000000000000",26492 => "0000000000000000",
26493 => "0000000000000000",26494 => "0000000000000000",
26495 => "0000000000000000",26496 => "0000000000000000",
26497 => "0000000000000000",26498 => "0000000000000000",
26499 => "0000000000000000",26500 => "0000000000000000",
26501 => "0000000000000000",26502 => "0000000000000000",
26503 => "0000000000000000",26504 => "0000000000000000",
26505 => "0000000000000000",26506 => "0000000000000000",
26507 => "0000000000000000",26508 => "0000000000000000",
26509 => "0000000000000000",26510 => "0000000000000000",
26511 => "0000000000000000",26512 => "0000000000000000",
26513 => "0000000000000000",26514 => "0000000000000000",
26515 => "0000000000000000",26516 => "0000000000000000",
26517 => "0000000000000000",26518 => "0000000000000000",
26519 => "0000000000000000",26520 => "0000000000000000",
26521 => "0000000000000000",26522 => "0000000000000000",
26523 => "0000000000000000",26524 => "0000000000000000",
26525 => "0000000000000000",26526 => "0000000000000000",
26527 => "0000000000000000",26528 => "0000000000000000",
26529 => "0000000000000000",26530 => "0000000000000000",
26531 => "0000000000000000",26532 => "0000000000000000",
26533 => "0000000000000000",26534 => "0000000000000000",
26535 => "0000000000000000",26536 => "0000000000000000",
26537 => "0000000000000000",26538 => "0000000000000000",
26539 => "0000000000000000",26540 => "0000000000000000",
26541 => "0000000000000000",26542 => "0000000000000000",
26543 => "0000000000000000",26544 => "0000000000000000",
26545 => "0000000000000000",26546 => "0000000000000000",
26547 => "0000000000000000",26548 => "0000000000000000",
26549 => "0000000000000000",26550 => "0000000000000000",
26551 => "0000000000000000",26552 => "0000000000000000",
26553 => "0000000000000000",26554 => "0000000000000000",
26555 => "0000000000000000",26556 => "0000000000000000",
26557 => "0000000000000000",26558 => "0000000000000000",
26559 => "0000000000000000",26560 => "0000000000000000",
26561 => "0000000000000000",26562 => "0000000000000000",
26563 => "0000000000000000",26564 => "0000000000000000",
26565 => "0000000000000000",26566 => "0000000000000000",
26567 => "0000000000000000",26568 => "0000000000000000",
26569 => "0000000000000000",26570 => "0000000000000000",
26571 => "0000000000000000",26572 => "0000000000000000",
26573 => "0000000000000000",26574 => "0000000000000000",
26575 => "0000000000000000",26576 => "0000000000000000",
26577 => "0000000000000000",26578 => "0000000000000000",
26579 => "0000000000000000",26580 => "0000000000000000",
26581 => "0000000000000000",26582 => "0000000000000000",
26583 => "0000000000000000",26584 => "0000000000000000",
26585 => "0000000000000000",26586 => "0000000000000000",
26587 => "0000000000000000",26588 => "0000000000000000",
26589 => "0000000000000000",26590 => "0000000000000000",
26591 => "0000000000000000",26592 => "0000000000000000",
26593 => "0000000000000000",26594 => "0000000000000000",
26595 => "0000000000000000",26596 => "0000000000000000",
26597 => "0000000000000000",26598 => "0000000000000000",
26599 => "0000000000000000",26600 => "0000000000000000",
26601 => "0000000000000000",26602 => "0000000000000000",
26603 => "0000000000000000",26604 => "0000000000000000",
26605 => "0000000000000000",26606 => "0000000000000000",
26607 => "0000000000000000",26608 => "0000000000000000",
26609 => "0000000000000000",26610 => "0000000000000000",
26611 => "0000000000000000",26612 => "0000000000000000",
26613 => "0000000000000000",26614 => "0000000000000000",
26615 => "0000000000000000",26616 => "0000000000000000",
26617 => "0000000000000000",26618 => "0000000000000000",
26619 => "0000000000000000",26620 => "0000000000000000",
26621 => "0000000000000000",26622 => "0000000000000000",
26623 => "0000000000000000",26624 => "0000000000000000",
26625 => "0000000000000000",26626 => "0000000000000000",
26627 => "0000000000000000",26628 => "0000000000000000",
26629 => "0000000000000000",26630 => "0000000000000000",
26631 => "0000000000000000",26632 => "0000000000000000",
26633 => "0000000000000000",26634 => "0000000000000000",
26635 => "0000000000000000",26636 => "0000000000000000",
26637 => "0000000000000000",26638 => "0000000000000000",
26639 => "0000000000000000",26640 => "0000000000000000",
26641 => "0000000000000000",26642 => "0000000000000000",
26643 => "0000000000000000",26644 => "0000000000000000",
26645 => "0000000000000000",26646 => "0000000000000000",
26647 => "0000000000000000",26648 => "0000000000000000",
26649 => "0000000000000000",26650 => "0000000000000000",
26651 => "0000000000000000",26652 => "0000000000000000",
26653 => "0000000000000000",26654 => "0000000000000000",
26655 => "0000000000000000",26656 => "0000000000000000",
26657 => "0000000000000000",26658 => "0000000000000000",
26659 => "0000000000000000",26660 => "0000000000000000",
26661 => "0000000000000000",26662 => "0000000000000000",
26663 => "0000000000000000",26664 => "0000000000000000",
26665 => "0000000000000000",26666 => "0000000000000000",
26667 => "0000000000000000",26668 => "0000000000000000",
26669 => "0000000000000000",26670 => "0000000000000000",
26671 => "0000000000000000",26672 => "0000000000000000",
26673 => "0000000000000000",26674 => "0000000000000000",
26675 => "0000000000000000",26676 => "0000000000000000",
26677 => "0000000000000000",26678 => "0000000000000000",
26679 => "0000000000000000",26680 => "0000000000000000",
26681 => "0000000000000000",26682 => "0000000000000000",
26683 => "0000000000000000",26684 => "0000000000000000",
26685 => "0000000000000000",26686 => "0000000000000000",
26687 => "0000000000000000",26688 => "0000000000000000",
26689 => "0000000000000000",26690 => "0000000000000000",
26691 => "0000000000000000",26692 => "0000000000000000",
26693 => "0000000000000000",26694 => "0000000000000000",
26695 => "0000000000000000",26696 => "0000000000000000",
26697 => "0000000000000000",26698 => "0000000000000000",
26699 => "0000000000000000",26700 => "0000000000000000",
26701 => "0000000000000000",26702 => "0000000000000000",
26703 => "0000000000000000",26704 => "0000000000000000",
26705 => "0000000000000000",26706 => "0000000000000000",
26707 => "0000000000000000",26708 => "0000000000000000",
26709 => "0000000000000000",26710 => "0000000000000000",
26711 => "0000000000000000",26712 => "0000000000000000",
26713 => "0000000000000000",26714 => "0000000000000000",
26715 => "0000000000000000",26716 => "0000000000000000",
26717 => "0000000000000000",26718 => "0000000000000000",
26719 => "0000000000000000",26720 => "0000000000000000",
26721 => "0000000000000000",26722 => "0000000000000000",
26723 => "0000000000000000",26724 => "0000000000000000",
26725 => "0000000000000000",26726 => "0000000000000000",
26727 => "0000000000000000",26728 => "0000000000000000",
26729 => "0000000000000000",26730 => "0000000000000000",
26731 => "0000000000000000",26732 => "0000000000000000",
26733 => "0000000000000000",26734 => "0000000000000000",
26735 => "0000000000000000",26736 => "0000000000000000",
26737 => "0000000000000000",26738 => "0000000000000000",
26739 => "0000000000000000",26740 => "0000000000000000",
26741 => "0000000000000000",26742 => "0000000000000000",
26743 => "0000000000000000",26744 => "0000000000000000",
26745 => "0000000000000000",26746 => "0000000000000000",
26747 => "0000000000000000",26748 => "0000000000000000",
26749 => "0000000000000000",26750 => "0000000000000000",
26751 => "0000000000000000",26752 => "0000000000000000",
26753 => "0000000000000000",26754 => "0000000000000000",
26755 => "0000000000000000",26756 => "0000000000000000",
26757 => "0000000000000000",26758 => "0000000000000000",
26759 => "0000000000000000",26760 => "0000000000000000",
26761 => "0000000000000000",26762 => "0000000000000000",
26763 => "0000000000000000",26764 => "0000000000000000",
26765 => "0000000000000000",26766 => "0000000000000000",
26767 => "0000000000000000",26768 => "0000000000000000",
26769 => "0000000000000000",26770 => "0000000000000000",
26771 => "0000000000000000",26772 => "0000000000000000",
26773 => "0000000000000000",26774 => "0000000000000000",
26775 => "0000000000000000",26776 => "0000000000000000",
26777 => "0000000000000000",26778 => "0000000000000000",
26779 => "0000000000000000",26780 => "0000000000000000",
26781 => "0000000000000000",26782 => "0000000000000000",
26783 => "0000000000000000",26784 => "0000000000000000",
26785 => "0000000000000000",26786 => "0000000000000000",
26787 => "0000000000000000",26788 => "0000000000000000",
26789 => "0000000000000000",26790 => "0000000000000000",
26791 => "0000000000000000",26792 => "0000000000000000",
26793 => "0000000000000000",26794 => "0000000000000000",
26795 => "0000000000000000",26796 => "0000000000000000",
26797 => "0000000000000000",26798 => "0000000000000000",
26799 => "0000000000000000",26800 => "0000000000000000",
26801 => "0000000000000000",26802 => "0000000000000000",
26803 => "0000000000000000",26804 => "0000000000000000",
26805 => "0000000000000000",26806 => "0000000000000000",
26807 => "0000000000000000",26808 => "0000000000000000",
26809 => "0000000000000000",26810 => "0000000000000000",
26811 => "0000000000000000",26812 => "0000000000000000",
26813 => "0000000000000000",26814 => "0000000000000000",
26815 => "0000000000000000",26816 => "0000000000000000",
26817 => "0000000000000000",26818 => "0000000000000000",
26819 => "0000000000000000",26820 => "0000000000000000",
26821 => "0000000000000000",26822 => "0000000000000000",
26823 => "0000000000000000",26824 => "0000000000000000",
26825 => "0000000000000000",26826 => "0000000000000000",
26827 => "0000000000000000",26828 => "0000000000000000",
26829 => "0000000000000000",26830 => "0000000000000000",
26831 => "0000000000000000",26832 => "0000000000000000",
26833 => "0000000000000000",26834 => "0000000000000000",
26835 => "0000000000000000",26836 => "0000000000000000",
26837 => "0000000000000000",26838 => "0000000000000000",
26839 => "0000000000000000",26840 => "0000000000000000",
26841 => "0000000000000000",26842 => "0000000000000000",
26843 => "0000000000000000",26844 => "0000000000000000",
26845 => "0000000000000000",26846 => "0000000000000000",
26847 => "0000000000000000",26848 => "0000000000000000",
26849 => "0000000000000000",26850 => "0000000000000000",
26851 => "0000000000000000",26852 => "0000000000000000",
26853 => "0000000000000000",26854 => "0000000000000000",
26855 => "0000000000000000",26856 => "0000000000000000",
26857 => "0000000000000000",26858 => "0000000000000000",
26859 => "0000000000000000",26860 => "0000000000000000",
26861 => "0000000000000000",26862 => "0000000000000000",
26863 => "0000000000000000",26864 => "0000000000000000",
26865 => "0000000000000000",26866 => "0000000000000000",
26867 => "0000000000000000",26868 => "0000000000000000",
26869 => "0000000000000000",26870 => "0000000000000000",
26871 => "0000000000000000",26872 => "0000000000000000",
26873 => "0000000000000000",26874 => "0000000000000000",
26875 => "0000000000000000",26876 => "0000000000000000",
26877 => "0000000000000000",26878 => "0000000000000000",
26879 => "0000000000000000",26880 => "0000000000000000",
26881 => "0000000000000000",26882 => "0000000000000000",
26883 => "0000000000000000",26884 => "0000000000000000",
26885 => "0000000000000000",26886 => "0000000000000000",
26887 => "0000000000000000",26888 => "0000000000000000",
26889 => "0000000000000000",26890 => "0000000000000000",
26891 => "0000000000000000",26892 => "0000000000000000",
26893 => "0000000000000000",26894 => "0000000000000000",
26895 => "0000000000000000",26896 => "0000000000000000",
26897 => "0000000000000000",26898 => "0000000000000000",
26899 => "0000000000000000",26900 => "0000000000000000",
26901 => "0000000000000000",26902 => "0000000000000000",
26903 => "0000000000000000",26904 => "0000000000000000",
26905 => "0000000000000000",26906 => "0000000000000000",
26907 => "0000000000000000",26908 => "0000000000000000",
26909 => "0000000000000000",26910 => "0000000000000000",
26911 => "0000000000000000",26912 => "0000000000000000",
26913 => "0000000000000000",26914 => "0000000000000000",
26915 => "0000000000000000",26916 => "0000000000000000",
26917 => "0000000000000000",26918 => "0000000000000000",
26919 => "0000000000000000",26920 => "0000000000000000",
26921 => "0000000000000000",26922 => "0000000000000000",
26923 => "0000000000000000",26924 => "0000000000000000",
26925 => "0000000000000000",26926 => "0000000000000000",
26927 => "0000000000000000",26928 => "0000000000000000",
26929 => "0000000000000000",26930 => "0000000000000000",
26931 => "0000000000000000",26932 => "0000000000000000",
26933 => "0000000000000000",26934 => "0000000000000000",
26935 => "0000000000000000",26936 => "0000000000000000",
26937 => "0000000000000000",26938 => "0000000000000000",
26939 => "0000000000000000",26940 => "0000000000000000",
26941 => "0000000000000000",26942 => "0000000000000000",
26943 => "0000000000000000",26944 => "0000000000000000",
26945 => "0000000000000000",26946 => "0000000000000000",
26947 => "0000000000000000",26948 => "0000000000000000",
26949 => "0000000000000000",26950 => "0000000000000000",
26951 => "0000000000000000",26952 => "0000000000000000",
26953 => "0000000000000000",26954 => "0000000000000000",
26955 => "0000000000000000",26956 => "0000000000000000",
26957 => "0000000000000000",26958 => "0000000000000000",
26959 => "0000000000000000",26960 => "0000000000000000",
26961 => "0000000000000000",26962 => "0000000000000000",
26963 => "0000000000000000",26964 => "0000000000000000",
26965 => "0000000000000000",26966 => "0000000000000000",
26967 => "0000000000000000",26968 => "0000000000000000",
26969 => "0000000000000000",26970 => "0000000000000000",
26971 => "0000000000000000",26972 => "0000000000000000",
26973 => "0000000000000000",26974 => "0000000000000000",
26975 => "0000000000000000",26976 => "0000000000000000",
26977 => "0000000000000000",26978 => "0000000000000000",
26979 => "0000000000000000",26980 => "0000000000000000",
26981 => "0000000000000000",26982 => "0000000000000000",
26983 => "0000000000000000",26984 => "0000000000000000",
26985 => "0000000000000000",26986 => "0000000000000000",
26987 => "0000000000000000",26988 => "0000000000000000",
26989 => "0000000000000000",26990 => "0000000000000000",
26991 => "0000000000000000",26992 => "0000000000000000",
26993 => "0000000000000000",26994 => "0000000000000000",
26995 => "0000000000000000",26996 => "0000000000000000",
26997 => "0000000000000000",26998 => "0000000000000000",
26999 => "0000000000000000",27000 => "0000000000000000",
27001 => "0000000000000000",27002 => "0000000000000000",
27003 => "0000000000000000",27004 => "0000000000000000",
27005 => "0000000000000000",27006 => "0000000000000000",
27007 => "0000000000000000",27008 => "0000000000000000",
27009 => "0000000000000000",27010 => "0000000000000000",
27011 => "0000000000000000",27012 => "0000000000000000",
27013 => "0000000000000000",27014 => "0000000000000000",
27015 => "0000000000000000",27016 => "0000000000000000",
27017 => "0000000000000000",27018 => "0000000000000000",
27019 => "0000000000000000",27020 => "0000000000000000",
27021 => "0000000000000000",27022 => "0000000000000000",
27023 => "0000000000000000",27024 => "0000000000000000",
27025 => "0000000000000000",27026 => "0000000000000000",
27027 => "0000000000000000",27028 => "0000000000000000",
27029 => "0000000000000000",27030 => "0000000000000000",
27031 => "0000000000000000",27032 => "0000000000000000",
27033 => "0000000000000000",27034 => "0000000000000000",
27035 => "0000000000000000",27036 => "0000000000000000",
27037 => "0000000000000000",27038 => "0000000000000000",
27039 => "0000000000000000",27040 => "0000000000000000",
27041 => "0000000000000000",27042 => "0000000000000000",
27043 => "0000000000000000",27044 => "0000000000000000",
27045 => "0000000000000000",27046 => "0000000000000000",
27047 => "0000000000000000",27048 => "0000000000000000",
27049 => "0000000000000000",27050 => "0000000000000000",
27051 => "0000000000000000",27052 => "0000000000000000",
27053 => "0000000000000000",27054 => "0000000000000000",
27055 => "0000000000000000",27056 => "0000000000000000",
27057 => "0000000000000000",27058 => "0000000000000000",
27059 => "0000000000000000",27060 => "0000000000000000",
27061 => "0000000000000000",27062 => "0000000000000000",
27063 => "0000000000000000",27064 => "0000000000000000",
27065 => "0000000000000000",27066 => "0000000000000000",
27067 => "0000000000000000",27068 => "0000000000000000",
27069 => "0000000000000000",27070 => "0000000000000000",
27071 => "0000000000000000",27072 => "0000000000000000",
27073 => "0000000000000000",27074 => "0000000000000000",
27075 => "0000000000000000",27076 => "0000000000000000",
27077 => "0000000000000000",27078 => "0000000000000000",
27079 => "0000000000000000",27080 => "0000000000000000",
27081 => "0000000000000000",27082 => "0000000000000000",
27083 => "0000000000000000",27084 => "0000000000000000",
27085 => "0000000000000000",27086 => "0000000000000000",
27087 => "0000000000000000",27088 => "0000000000000000",
27089 => "0000000000000000",27090 => "0000000000000000",
27091 => "0000000000000000",27092 => "0000000000000000",
27093 => "0000000000000000",27094 => "0000000000000000",
27095 => "0000000000000000",27096 => "0000000000000000",
27097 => "0000000000000000",27098 => "0000000000000000",
27099 => "0000000000000000",27100 => "0000000000000000",
27101 => "0000000000000000",27102 => "0000000000000000",
27103 => "0000000000000000",27104 => "0000000000000000",
27105 => "0000000000000000",27106 => "0000000000000000",
27107 => "0000000000000000",27108 => "0000000000000000",
27109 => "0000000000000000",27110 => "0000000000000000",
27111 => "0000000000000000",27112 => "0000000000000000",
27113 => "0000000000000000",27114 => "0000000000000000",
27115 => "0000000000000000",27116 => "0000000000000000",
27117 => "0000000000000000",27118 => "0000000000000000",
27119 => "0000000000000000",27120 => "0000000000000000",
27121 => "0000000000000000",27122 => "0000000000000000",
27123 => "0000000000000000",27124 => "0000000000000000",
27125 => "0000000000000000",27126 => "0000000000000000",
27127 => "0000000000000000",27128 => "0000000000000000",
27129 => "0000000000000000",27130 => "0000000000000000",
27131 => "0000000000000000",27132 => "0000000000000000",
27133 => "0000000000000000",27134 => "0000000000000000",
27135 => "0000000000000000",27136 => "0000000000000000",
27137 => "0000000000000000",27138 => "0000000000000000",
27139 => "0000000000000000",27140 => "0000000000000000",
27141 => "0000000000000000",27142 => "0000000000000000",
27143 => "0000000000000000",27144 => "0000000000000000",
27145 => "0000000000000000",27146 => "0000000000000000",
27147 => "0000000000000000",27148 => "0000000000000000",
27149 => "0000000000000000",27150 => "0000000000000000",
27151 => "0000000000000000",27152 => "0000000000000000",
27153 => "0000000000000000",27154 => "0000000000000000",
27155 => "0000000000000000",27156 => "0000000000000000",
27157 => "0000000000000000",27158 => "0000000000000000",
27159 => "0000000000000000",27160 => "0000000000000000",
27161 => "0000000000000000",27162 => "0000000000000000",
27163 => "0000000000000000",27164 => "0000000000000000",
27165 => "0000000000000000",27166 => "0000000000000000",
27167 => "0000000000000000",27168 => "0000000000000000",
27169 => "0000000000000000",27170 => "0000000000000000",
27171 => "0000000000000000",27172 => "0000000000000000",
27173 => "0000000000000000",27174 => "0000000000000000",
27175 => "0000000000000000",27176 => "0000000000000000",
27177 => "0000000000000000",27178 => "0000000000000000",
27179 => "0000000000000000",27180 => "0000000000000000",
27181 => "0000000000000000",27182 => "0000000000000000",
27183 => "0000000000000000",27184 => "0000000000000000",
27185 => "0000000000000000",27186 => "0000000000000000",
27187 => "0000000000000000",27188 => "0000000000000000",
27189 => "0000000000000000",27190 => "0000000000000000",
27191 => "0000000000000000",27192 => "0000000000000000",
27193 => "0000000000000000",27194 => "0000000000000000",
27195 => "0000000000000000",27196 => "0000000000000000",
27197 => "0000000000000000",27198 => "0000000000000000",
27199 => "0000000000000000",27200 => "0000000000000000",
27201 => "0000000000000000",27202 => "0000000000000000",
27203 => "0000000000000000",27204 => "0000000000000000",
27205 => "0000000000000000",27206 => "0000000000000000",
27207 => "0000000000000000",27208 => "0000000000000000",
27209 => "0000000000000000",27210 => "0000000000000000",
27211 => "0000000000000000",27212 => "0000000000000000",
27213 => "0000000000000000",27214 => "0000000000000000",
27215 => "0000000000000000",27216 => "0000000000000000",
27217 => "0000000000000000",27218 => "0000000000000000",
27219 => "0000000000000000",27220 => "0000000000000000",
27221 => "0000000000000000",27222 => "0000000000000000",
27223 => "0000000000000000",27224 => "0000000000000000",
27225 => "0000000000000000",27226 => "0000000000000000",
27227 => "0000000000000000",27228 => "0000000000000000",
27229 => "0000000000000000",27230 => "0000000000000000",
27231 => "0000000000000000",27232 => "0000000000000000",
27233 => "0000000000000000",27234 => "0000000000000000",
27235 => "0000000000000000",27236 => "0000000000000000",
27237 => "0000000000000000",27238 => "0000000000000000",
27239 => "0000000000000000",27240 => "0000000000000000",
27241 => "0000000000000000",27242 => "0000000000000000",
27243 => "0000000000000000",27244 => "0000000000000000",
27245 => "0000000000000000",27246 => "0000000000000000",
27247 => "0000000000000000",27248 => "0000000000000000",
27249 => "0000000000000000",27250 => "0000000000000000",
27251 => "0000000000000000",27252 => "0000000000000000",
27253 => "0000000000000000",27254 => "0000000000000000",
27255 => "0000000000000000",27256 => "0000000000000000",
27257 => "0000000000000000",27258 => "0000000000000000",
27259 => "0000000000000000",27260 => "0000000000000000",
27261 => "0000000000000000",27262 => "0000000000000000",
27263 => "0000000000000000",27264 => "0000000000000000",
27265 => "0000000000000000",27266 => "0000000000000000",
27267 => "0000000000000000",27268 => "0000000000000000",
27269 => "0000000000000000",27270 => "0000000000000000",
27271 => "0000000000000000",27272 => "0000000000000000",
27273 => "0000000000000000",27274 => "0000000000000000",
27275 => "0000000000000000",27276 => "0000000000000000",
27277 => "0000000000000000",27278 => "0000000000000000",
27279 => "0000000000000000",27280 => "0000000000000000",
27281 => "0000000000000000",27282 => "0000000000000000",
27283 => "0000000000000000",27284 => "0000000000000000",
27285 => "0000000000000000",27286 => "0000000000000000",
27287 => "0000000000000000",27288 => "0000000000000000",
27289 => "0000000000000000",27290 => "0000000000000000",
27291 => "0000000000000000",27292 => "0000000000000000",
27293 => "0000000000000000",27294 => "0000000000000000",
27295 => "0000000000000000",27296 => "0000000000000000",
27297 => "0000000000000000",27298 => "0000000000000000",
27299 => "0000000000000000",27300 => "0000000000000000",
27301 => "0000000000000000",27302 => "0000000000000000",
27303 => "0000000000000000",27304 => "0000000000000000",
27305 => "0000000000000000",27306 => "0000000000000000",
27307 => "0000000000000000",27308 => "0000000000000000",
27309 => "0000000000000000",27310 => "0000000000000000",
27311 => "0000000000000000",27312 => "0000000000000000",
27313 => "0000000000000000",27314 => "0000000000000000",
27315 => "0000000000000000",27316 => "0000000000000000",
27317 => "0000000000000000",27318 => "0000000000000000",
27319 => "0000000000000000",27320 => "0000000000000000",
27321 => "0000000000000000",27322 => "0000000000000000",
27323 => "0000000000000000",27324 => "0000000000000000",
27325 => "0000000000000000",27326 => "0000000000000000",
27327 => "0000000000000000",27328 => "0000000000000000",
27329 => "0000000000000000",27330 => "0000000000000000",
27331 => "0000000000000000",27332 => "0000000000000000",
27333 => "0000000000000000",27334 => "0000000000000000",
27335 => "0000000000000000",27336 => "0000000000000000",
27337 => "0000000000000000",27338 => "0000000000000000",
27339 => "0000000000000000",27340 => "0000000000000000",
27341 => "0000000000000000",27342 => "0000000000000000",
27343 => "0000000000000000",27344 => "0000000000000000",
27345 => "0000000000000000",27346 => "0000000000000000",
27347 => "0000000000000000",27348 => "0000000000000000",
27349 => "0000000000000000",27350 => "0000000000000000",
27351 => "0000000000000000",27352 => "0000000000000000",
27353 => "0000000000000000",27354 => "0000000000000000",
27355 => "0000000000000000",27356 => "0000000000000000",
27357 => "0000000000000000",27358 => "0000000000000000",
27359 => "0000000000000000",27360 => "0000000000000000",
27361 => "0000000000000000",27362 => "0000000000000000",
27363 => "0000000000000000",27364 => "0000000000000000",
27365 => "0000000000000000",27366 => "0000000000000000",
27367 => "0000000000000000",27368 => "0000000000000000",
27369 => "0000000000000000",27370 => "0000000000000000",
27371 => "0000000000000000",27372 => "0000000000000000",
27373 => "0000000000000000",27374 => "0000000000000000",
27375 => "0000000000000000",27376 => "0000000000000000",
27377 => "0000000000000000",27378 => "0000000000000000",
27379 => "0000000000000000",27380 => "0000000000000000",
27381 => "0000000000000000",27382 => "0000000000000000",
27383 => "0000000000000000",27384 => "0000000000000000",
27385 => "0000000000000000",27386 => "0000000000000000",
27387 => "0000000000000000",27388 => "0000000000000000",
27389 => "0000000000000000",27390 => "0000000000000000",
27391 => "0000000000000000",27392 => "0000000000000000",
27393 => "0000000000000000",27394 => "0000000000000000",
27395 => "0000000000000000",27396 => "0000000000000000",
27397 => "0000000000000000",27398 => "0000000000000000",
27399 => "0000000000000000",27400 => "0000000000000000",
27401 => "0000000000000000",27402 => "0000000000000000",
27403 => "0000000000000000",27404 => "0000000000000000",
27405 => "0000000000000000",27406 => "0000000000000000",
27407 => "0000000000000000",27408 => "0000000000000000",
27409 => "0000000000000000",27410 => "0000000000000000",
27411 => "0000000000000000",27412 => "0000000000000000",
27413 => "0000000000000000",27414 => "0000000000000000",
27415 => "0000000000000000",27416 => "0000000000000000",
27417 => "0000000000000000",27418 => "0000000000000000",
27419 => "0000000000000000",27420 => "0000000000000000",
27421 => "0000000000000000",27422 => "0000000000000000",
27423 => "0000000000000000",27424 => "0000000000000000",
27425 => "0000000000000000",27426 => "0000000000000000",
27427 => "0000000000000000",27428 => "0000000000000000",
27429 => "0000000000000000",27430 => "0000000000000000",
27431 => "0000000000000000",27432 => "0000000000000000",
27433 => "0000000000000000",27434 => "0000000000000000",
27435 => "0000000000000000",27436 => "0000000000000000",
27437 => "0000000000000000",27438 => "0000000000000000",
27439 => "0000000000000000",27440 => "0000000000000000",
27441 => "0000000000000000",27442 => "0000000000000000",
27443 => "0000000000000000",27444 => "0000000000000000",
27445 => "0000000000000000",27446 => "0000000000000000",
27447 => "0000000000000000",27448 => "0000000000000000",
27449 => "0000000000000000",27450 => "0000000000000000",
27451 => "0000000000000000",27452 => "0000000000000000",
27453 => "0000000000000000",27454 => "0000000000000000",
27455 => "0000000000000000",27456 => "0000000000000000",
27457 => "0000000000000000",27458 => "0000000000000000",
27459 => "0000000000000000",27460 => "0000000000000000",
27461 => "0000000000000000",27462 => "0000000000000000",
27463 => "0000000000000000",27464 => "0000000000000000",
27465 => "0000000000000000",27466 => "0000000000000000",
27467 => "0000000000000000",27468 => "0000000000000000",
27469 => "0000000000000000",27470 => "0000000000000000",
27471 => "0000000000000000",27472 => "0000000000000000",
27473 => "0000000000000000",27474 => "0000000000000000",
27475 => "0000000000000000",27476 => "0000000000000000",
27477 => "0000000000000000",27478 => "0000000000000000",
27479 => "0000000000000000",27480 => "0000000000000000",
27481 => "0000000000000000",27482 => "0000000000000000",
27483 => "0000000000000000",27484 => "0000000000000000",
27485 => "0000000000000000",27486 => "0000000000000000",
27487 => "0000000000000000",27488 => "0000000000000000",
27489 => "0000000000000000",27490 => "0000000000000000",
27491 => "0000000000000000",27492 => "0000000000000000",
27493 => "0000000000000000",27494 => "0000000000000000",
27495 => "0000000000000000",27496 => "0000000000000000",
27497 => "0000000000000000",27498 => "0000000000000000",
27499 => "0000000000000000",27500 => "0000000000000000",
27501 => "0000000000000000",27502 => "0000000000000000",
27503 => "0000000000000000",27504 => "0000000000000000",
27505 => "0000000000000000",27506 => "0000000000000000",
27507 => "0000000000000000",27508 => "0000000000000000",
27509 => "0000000000000000",27510 => "0000000000000000",
27511 => "0000000000000000",27512 => "0000000000000000",
27513 => "0000000000000000",27514 => "0000000000000000",
27515 => "0000000000000000",27516 => "0000000000000000",
27517 => "0000000000000000",27518 => "0000000000000000",
27519 => "0000000000000000",27520 => "0000000000000000",
27521 => "0000000000000000",27522 => "0000000000000000",
27523 => "0000000000000000",27524 => "0000000000000000",
27525 => "0000000000000000",27526 => "0000000000000000",
27527 => "0000000000000000",27528 => "0000000000000000",
27529 => "0000000000000000",27530 => "0000000000000000",
27531 => "0000000000000000",27532 => "0000000000000000",
27533 => "0000000000000000",27534 => "0000000000000000",
27535 => "0000000000000000",27536 => "0000000000000000",
27537 => "0000000000000000",27538 => "0000000000000000",
27539 => "0000000000000000",27540 => "0000000000000000",
27541 => "0000000000000000",27542 => "0000000000000000",
27543 => "0000000000000000",27544 => "0000000000000000",
27545 => "0000000000000000",27546 => "0000000000000000",
27547 => "0000000000000000",27548 => "0000000000000000",
27549 => "0000000000000000",27550 => "0000000000000000",
27551 => "0000000000000000",27552 => "0000000000000000",
27553 => "0000000000000000",27554 => "0000000000000000",
27555 => "0000000000000000",27556 => "0000000000000000",
27557 => "0000000000000000",27558 => "0000000000000000",
27559 => "0000000000000000",27560 => "0000000000000000",
27561 => "0000000000000000",27562 => "0000000000000000",
27563 => "0000000000000000",27564 => "0000000000000000",
27565 => "0000000000000000",27566 => "0000000000000000",
27567 => "0000000000000000",27568 => "0000000000000000",
27569 => "0000000000000000",27570 => "0000000000000000",
27571 => "0000000000000000",27572 => "0000000000000000",
27573 => "0000000000000000",27574 => "0000000000000000",
27575 => "0000000000000000",27576 => "0000000000000000",
27577 => "0000000000000000",27578 => "0000000000000000",
27579 => "0000000000000000",27580 => "0000000000000000",
27581 => "0000000000000000",27582 => "0000000000000000",
27583 => "0000000000000000",27584 => "0000000000000000",
27585 => "0000000000000000",27586 => "0000000000000000",
27587 => "0000000000000000",27588 => "0000000000000000",
27589 => "0000000000000000",27590 => "0000000000000000",
27591 => "0000000000000000",27592 => "0000000000000000",
27593 => "0000000000000000",27594 => "0000000000000000",
27595 => "0000000000000000",27596 => "0000000000000000",
27597 => "0000000000000000",27598 => "0000000000000000",
27599 => "0000000000000000",27600 => "0000000000000000",
27601 => "0000000000000000",27602 => "0000000000000000",
27603 => "0000000000000000",27604 => "0000000000000000",
27605 => "0000000000000000",27606 => "0000000000000000",
27607 => "0000000000000000",27608 => "0000000000000000",
27609 => "0000000000000000",27610 => "0000000000000000",
27611 => "0000000000000000",27612 => "0000000000000000",
27613 => "0000000000000000",27614 => "0000000000000000",
27615 => "0000000000000000",27616 => "0000000000000000",
27617 => "0000000000000000",27618 => "0000000000000000",
27619 => "0000000000000000",27620 => "0000000000000000",
27621 => "0000000000000000",27622 => "0000000000000000",
27623 => "0000000000000000",27624 => "0000000000000000",
27625 => "0000000000000000",27626 => "0000000000000000",
27627 => "0000000000000000",27628 => "0000000000000000",
27629 => "0000000000000000",27630 => "0000000000000000",
27631 => "0000000000000000",27632 => "0000000000000000",
27633 => "0000000000000000",27634 => "0000000000000000",
27635 => "0000000000000000",27636 => "0000000000000000",
27637 => "0000000000000000",27638 => "0000000000000000",
27639 => "0000000000000000",27640 => "0000000000000000",
27641 => "0000000000000000",27642 => "0000000000000000",
27643 => "0000000000000000",27644 => "0000000000000000",
27645 => "0000000000000000",27646 => "0000000000000000",
27647 => "0000000000000000",27648 => "0000000000000000",
27649 => "0000000000000000",27650 => "0000000000000000",
27651 => "0000000000000000",27652 => "0000000000000000",
27653 => "0000000000000000",27654 => "0000000000000000",
27655 => "0000000000000000",27656 => "0000000000000000",
27657 => "0000000000000000",27658 => "0000000000000000",
27659 => "0000000000000000",27660 => "0000000000000000",
27661 => "0000000000000000",27662 => "0000000000000000",
27663 => "0000000000000000",27664 => "0000000000000000",
27665 => "0000000000000000",27666 => "0000000000000000",
27667 => "0000000000000000",27668 => "0000000000000000",
27669 => "0000000000000000",27670 => "0000000000000000",
27671 => "0000000000000000",27672 => "0000000000000000",
27673 => "0000000000000000",27674 => "0000000000000000",
27675 => "0000000000000000",27676 => "0000000000000000",
27677 => "0000000000000000",27678 => "0000000000000000",
27679 => "0000000000000000",27680 => "0000000000000000",
27681 => "0000000000000000",27682 => "0000000000000000",
27683 => "0000000000000000",27684 => "0000000000000000",
27685 => "0000000000000000",27686 => "0000000000000000",
27687 => "0000000000000000",27688 => "0000000000000000",
27689 => "0000000000000000",27690 => "0000000000000000",
27691 => "0000000000000000",27692 => "0000000000000000",
27693 => "0000000000000000",27694 => "0000000000000000",
27695 => "0000000000000000",27696 => "0000000000000000",
27697 => "0000000000000000",27698 => "0000000000000000",
27699 => "0000000000000000",27700 => "0000000000000000",
27701 => "0000000000000000",27702 => "0000000000000000",
27703 => "0000000000000000",27704 => "0000000000000000",
27705 => "0000000000000000",27706 => "0000000000000000",
27707 => "0000000000000000",27708 => "0000000000000000",
27709 => "0000000000000000",27710 => "0000000000000000",
27711 => "0000000000000000",27712 => "0000000000000000",
27713 => "0000000000000000",27714 => "0000000000000000",
27715 => "0000000000000000",27716 => "0000000000000000",
27717 => "0000000000000000",27718 => "0000000000000000",
27719 => "0000000000000000",27720 => "0000000000000000",
27721 => "0000000000000000",27722 => "0000000000000000",
27723 => "0000000000000000",27724 => "0000000000000000",
27725 => "0000000000000000",27726 => "0000000000000000",
27727 => "0000000000000000",27728 => "0000000000000000",
27729 => "0000000000000000",27730 => "0000000000000000",
27731 => "0000000000000000",27732 => "0000000000000000",
27733 => "0000000000000000",27734 => "0000000000000000",
27735 => "0000000000000000",27736 => "0000000000000000",
27737 => "0000000000000000",27738 => "0000000000000000",
27739 => "0000000000000000",27740 => "0000000000000000",
27741 => "0000000000000000",27742 => "0000000000000000",
27743 => "0000000000000000",27744 => "0000000000000000",
27745 => "0000000000000000",27746 => "0000000000000000",
27747 => "0000000000000000",27748 => "0000000000000000",
27749 => "0000000000000000",27750 => "0000000000000000",
27751 => "0000000000000000",27752 => "0000000000000000",
27753 => "0000000000000000",27754 => "0000000000000000",
27755 => "0000000000000000",27756 => "0000000000000000",
27757 => "0000000000000000",27758 => "0000000000000000",
27759 => "0000000000000000",27760 => "0000000000000000",
27761 => "0000000000000000",27762 => "0000000000000000",
27763 => "0000000000000000",27764 => "0000000000000000",
27765 => "0000000000000000",27766 => "0000000000000000",
27767 => "0000000000000000",27768 => "0000000000000000",
27769 => "0000000000000000",27770 => "0000000000000000",
27771 => "0000000000000000",27772 => "0000000000000000",
27773 => "0000000000000000",27774 => "0000000000000000",
27775 => "0000000000000000",27776 => "0000000000000000",
27777 => "0000000000000000",27778 => "0000000000000000",
27779 => "0000000000000000",27780 => "0000000000000000",
27781 => "0000000000000000",27782 => "0000000000000000",
27783 => "0000000000000000",27784 => "0000000000000000",
27785 => "0000000000000000",27786 => "0000000000000000",
27787 => "0000000000000000",27788 => "0000000000000000",
27789 => "0000000000000000",27790 => "0000000000000000",
27791 => "0000000000000000",27792 => "0000000000000000",
27793 => "0000000000000000",27794 => "0000000000000000",
27795 => "0000000000000000",27796 => "0000000000000000",
27797 => "0000000000000000",27798 => "0000000000000000",
27799 => "0000000000000000",27800 => "0000000000000000",
27801 => "0000000000000000",27802 => "0000000000000000",
27803 => "0000000000000000",27804 => "0000000000000000",
27805 => "0000000000000000",27806 => "0000000000000000",
27807 => "0000000000000000",27808 => "0000000000000000",
27809 => "0000000000000000",27810 => "0000000000000000",
27811 => "0000000000000000",27812 => "0000000000000000",
27813 => "0000000000000000",27814 => "0000000000000000",
27815 => "0000000000000000",27816 => "0000000000000000",
27817 => "0000000000000000",27818 => "0000000000000000",
27819 => "0000000000000000",27820 => "0000000000000000",
27821 => "0000000000000000",27822 => "0000000000000000",
27823 => "0000000000000000",27824 => "0000000000000000",
27825 => "0000000000000000",27826 => "0000000000000000",
27827 => "0000000000000000",27828 => "0000000000000000",
27829 => "0000000000000000",27830 => "0000000000000000",
27831 => "0000000000000000",27832 => "0000000000000000",
27833 => "0000000000000000",27834 => "0000000000000000",
27835 => "0000000000000000",27836 => "0000000000000000",
27837 => "0000000000000000",27838 => "0000000000000000",
27839 => "0000000000000000",27840 => "0000000000000000",
27841 => "0000000000000000",27842 => "0000000000000000",
27843 => "0000000000000000",27844 => "0000000000000000",
27845 => "0000000000000000",27846 => "0000000000000000",
27847 => "0000000000000000",27848 => "0000000000000000",
27849 => "0000000000000000",27850 => "0000000000000000",
27851 => "0000000000000000",27852 => "0000000000000000",
27853 => "0000000000000000",27854 => "0000000000000000",
27855 => "0000000000000000",27856 => "0000000000000000",
27857 => "0000000000000000",27858 => "0000000000000000",
27859 => "0000000000000000",27860 => "0000000000000000",
27861 => "0000000000000000",27862 => "0000000000000000",
27863 => "0000000000000000",27864 => "0000000000000000",
27865 => "0000000000000000",27866 => "0000000000000000",
27867 => "0000000000000000",27868 => "0000000000000000",
27869 => "0000000000000000",27870 => "0000000000000000",
27871 => "0000000000000000",27872 => "0000000000000000",
27873 => "0000000000000000",27874 => "0000000000000000",
27875 => "0000000000000000",27876 => "0000000000000000",
27877 => "0000000000000000",27878 => "0000000000000000",
27879 => "0000000000000000",27880 => "0000000000000000",
27881 => "0000000000000000",27882 => "0000000000000000",
27883 => "0000000000000000",27884 => "0000000000000000",
27885 => "0000000000000000",27886 => "0000000000000000",
27887 => "0000000000000000",27888 => "0000000000000000",
27889 => "0000000000000000",27890 => "0000000000000000",
27891 => "0000000000000000",27892 => "0000000000000000",
27893 => "0000000000000000",27894 => "0000000000000000",
27895 => "0000000000000000",27896 => "0000000000000000",
27897 => "0000000000000000",27898 => "0000000000000000",
27899 => "0000000000000000",27900 => "0000000000000000",
27901 => "0000000000000000",27902 => "0000000000000000",
27903 => "0000000000000000",27904 => "0000000000000000",
27905 => "0000000000000000",27906 => "0000000000000000",
27907 => "0000000000000000",27908 => "0000000000000000",
27909 => "0000000000000000",27910 => "0000000000000000",
27911 => "0000000000000000",27912 => "0000000000000000",
27913 => "0000000000000000",27914 => "0000000000000000",
27915 => "0000000000000000",27916 => "0000000000000000",
27917 => "0000000000000000",27918 => "0000000000000000",
27919 => "0000000000000000",27920 => "0000000000000000",
27921 => "0000000000000000",27922 => "0000000000000000",
27923 => "0000000000000000",27924 => "0000000000000000",
27925 => "0000000000000000",27926 => "0000000000000000",
27927 => "0000000000000000",27928 => "0000000000000000",
27929 => "0000000000000000",27930 => "0000000000000000",
27931 => "0000000000000000",27932 => "0000000000000000",
27933 => "0000000000000000",27934 => "0000000000000000",
27935 => "0000000000000000",27936 => "0000000000000000",
27937 => "0000000000000000",27938 => "0000000000000000",
27939 => "0000000000000000",27940 => "0000000000000000",
27941 => "0000000000000000",27942 => "0000000000000000",
27943 => "0000000000000000",27944 => "0000000000000000",
27945 => "0000000000000000",27946 => "0000000000000000",
27947 => "0000000000000000",27948 => "0000000000000000",
27949 => "0000000000000000",27950 => "0000000000000000",
27951 => "0000000000000000",27952 => "0000000000000000",
27953 => "0000000000000000",27954 => "0000000000000000",
27955 => "0000000000000000",27956 => "0000000000000000",
27957 => "0000000000000000",27958 => "0000000000000000",
27959 => "0000000000000000",27960 => "0000000000000000",
27961 => "0000000000000000",27962 => "0000000000000000",
27963 => "0000000000000000",27964 => "0000000000000000",
27965 => "0000000000000000",27966 => "0000000000000000",
27967 => "0000000000000000",27968 => "0000000000000000",
27969 => "0000000000000000",27970 => "0000000000000000",
27971 => "0000000000000000",27972 => "0000000000000000",
27973 => "0000000000000000",27974 => "0000000000000000",
27975 => "0000000000000000",27976 => "0000000000000000",
27977 => "0000000000000000",27978 => "0000000000000000",
27979 => "0000000000000000",27980 => "0000000000000000",
27981 => "0000000000000000",27982 => "0000000000000000",
27983 => "0000000000000000",27984 => "0000000000000000",
27985 => "0000000000000000",27986 => "0000000000000000",
27987 => "0000000000000000",27988 => "0000000000000000",
27989 => "0000000000000000",27990 => "0000000000000000",
27991 => "0000000000000000",27992 => "0000000000000000",
27993 => "0000000000000000",27994 => "0000000000000000",
27995 => "0000000000000000",27996 => "0000000000000000",
27997 => "0000000000000000",27998 => "0000000000000000",
27999 => "0000000000000000",28000 => "0000000000000000",
28001 => "0000000000000000",28002 => "0000000000000000",
28003 => "0000000000000000",28004 => "0000000000000000",
28005 => "0000000000000000",28006 => "0000000000000000",
28007 => "0000000000000000",28008 => "0000000000000000",
28009 => "0000000000000000",28010 => "0000000000000000",
28011 => "0000000000000000",28012 => "0000000000000000",
28013 => "0000000000000000",28014 => "0000000000000000",
28015 => "0000000000000000",28016 => "0000000000000000",
28017 => "0000000000000000",28018 => "0000000000000000",
28019 => "0000000000000000",28020 => "0000000000000000",
28021 => "0000000000000000",28022 => "0000000000000000",
28023 => "0000000000000000",28024 => "0000000000000000",
28025 => "0000000000000000",28026 => "0000000000000000",
28027 => "0000000000000000",28028 => "0000000000000000",
28029 => "0000000000000000",28030 => "0000000000000000",
28031 => "0000000000000000",28032 => "0000000000000000",
28033 => "0000000000000000",28034 => "0000000000000000",
28035 => "0000000000000000",28036 => "0000000000000000",
28037 => "0000000000000000",28038 => "0000000000000000",
28039 => "0000000000000000",28040 => "0000000000000000",
28041 => "0000000000000000",28042 => "0000000000000000",
28043 => "0000000000000000",28044 => "0000000000000000",
28045 => "0000000000000000",28046 => "0000000000000000",
28047 => "0000000000000000",28048 => "0000000000000000",
28049 => "0000000000000000",28050 => "0000000000000000",
28051 => "0000000000000000",28052 => "0000000000000000",
28053 => "0000000000000000",28054 => "0000000000000000",
28055 => "0000000000000000",28056 => "0000000000000000",
28057 => "0000000000000000",28058 => "0000000000000000",
28059 => "0000000000000000",28060 => "0000000000000000",
28061 => "0000000000000000",28062 => "0000000000000000",
28063 => "0000000000000000",28064 => "0000000000000000",
28065 => "0000000000000000",28066 => "0000000000000000",
28067 => "0000000000000000",28068 => "0000000000000000",
28069 => "0000000000000000",28070 => "0000000000000000",
28071 => "0000000000000000",28072 => "0000000000000000",
28073 => "0000000000000000",28074 => "0000000000000000",
28075 => "0000000000000000",28076 => "0000000000000000",
28077 => "0000000000000000",28078 => "0000000000000000",
28079 => "0000000000000000",28080 => "0000000000000000",
28081 => "0000000000000000",28082 => "0000000000000000",
28083 => "0000000000000000",28084 => "0000000000000000",
28085 => "0000000000000000",28086 => "0000000000000000",
28087 => "0000000000000000",28088 => "0000000000000000",
28089 => "0000000000000000",28090 => "0000000000000000",
28091 => "0000000000000000",28092 => "0000000000000000",
28093 => "0000000000000000",28094 => "0000000000000000",
28095 => "0000000000000000",28096 => "0000000000000000",
28097 => "0000000000000000",28098 => "0000000000000000",
28099 => "0000000000000000",28100 => "0000000000000000",
28101 => "0000000000000000",28102 => "0000000000000000",
28103 => "0000000000000000",28104 => "0000000000000000",
28105 => "0000000000000000",28106 => "0000000000000000",
28107 => "0000000000000000",28108 => "0000000000000000",
28109 => "0000000000000000",28110 => "0000000000000000",
28111 => "0000000000000000",28112 => "0000000000000000",
28113 => "0000000000000000",28114 => "0000000000000000",
28115 => "0000000000000000",28116 => "0000000000000000",
28117 => "0000000000000000",28118 => "0000000000000000",
28119 => "0000000000000000",28120 => "0000000000000000",
28121 => "0000000000000000",28122 => "0000000000000000",
28123 => "0000000000000000",28124 => "0000000000000000",
28125 => "0000000000000000",28126 => "0000000000000000",
28127 => "0000000000000000",28128 => "0000000000000000",
28129 => "0000000000000000",28130 => "0000000000000000",
28131 => "0000000000000000",28132 => "0000000000000000",
28133 => "0000000000000000",28134 => "0000000000000000",
28135 => "0000000000000000",28136 => "0000000000000000",
28137 => "0000000000000000",28138 => "0000000000000000",
28139 => "0000000000000000",28140 => "0000000000000000",
28141 => "0000000000000000",28142 => "0000000000000000",
28143 => "0000000000000000",28144 => "0000000000000000",
28145 => "0000000000000000",28146 => "0000000000000000",
28147 => "0000000000000000",28148 => "0000000000000000",
28149 => "0000000000000000",28150 => "0000000000000000",
28151 => "0000000000000000",28152 => "0000000000000000",
28153 => "0000000000000000",28154 => "0000000000000000",
28155 => "0000000000000000",28156 => "0000000000000000",
28157 => "0000000000000000",28158 => "0000000000000000",
28159 => "0000000000000000",28160 => "0000000000000000",
28161 => "0000000000000000",28162 => "0000000000000000",
28163 => "0000000000000000",28164 => "0000000000000000",
28165 => "0000000000000000",28166 => "0000000000000000",
28167 => "0000000000000000",28168 => "0000000000000000",
28169 => "0000000000000000",28170 => "0000000000000000",
28171 => "0000000000000000",28172 => "0000000000000000",
28173 => "0000000000000000",28174 => "0000000000000000",
28175 => "0000000000000000",28176 => "0000000000000000",
28177 => "0000000000000000",28178 => "0000000000000000",
28179 => "0000000000000000",28180 => "0000000000000000",
28181 => "0000000000000000",28182 => "0000000000000000",
28183 => "0000000000000000",28184 => "0000000000000000",
28185 => "0000000000000000",28186 => "0000000000000000",
28187 => "0000000000000000",28188 => "0000000000000000",
28189 => "0000000000000000",28190 => "0000000000000000",
28191 => "0000000000000000",28192 => "0000000000000000",
28193 => "0000000000000000",28194 => "0000000000000000",
28195 => "0000000000000000",28196 => "0000000000000000",
28197 => "0000000000000000",28198 => "0000000000000000",
28199 => "0000000000000000",28200 => "0000000000000000",
28201 => "0000000000000000",28202 => "0000000000000000",
28203 => "0000000000000000",28204 => "0000000000000000",
28205 => "0000000000000000",28206 => "0000000000000000",
28207 => "0000000000000000",28208 => "0000000000000000",
28209 => "0000000000000000",28210 => "0000000000000000",
28211 => "0000000000000000",28212 => "0000000000000000",
28213 => "0000000000000000",28214 => "0000000000000000",
28215 => "0000000000000000",28216 => "0000000000000000",
28217 => "0000000000000000",28218 => "0000000000000000",
28219 => "0000000000000000",28220 => "0000000000000000",
28221 => "0000000000000000",28222 => "0000000000000000",
28223 => "0000000000000000",28224 => "0000000000000000",
28225 => "0000000000000000",28226 => "0000000000000000",
28227 => "0000000000000000",28228 => "0000000000000000",
28229 => "0000000000000000",28230 => "0000000000000000",
28231 => "0000000000000000",28232 => "0000000000000000",
28233 => "0000000000000000",28234 => "0000000000000000",
28235 => "0000000000000000",28236 => "0000000000000000",
28237 => "0000000000000000",28238 => "0000000000000000",
28239 => "0000000000000000",28240 => "0000000000000000",
28241 => "0000000000000000",28242 => "0000000000000000",
28243 => "0000000000000000",28244 => "0000000000000000",
28245 => "0000000000000000",28246 => "0000000000000000",
28247 => "0000000000000000",28248 => "0000000000000000",
28249 => "0000000000000000",28250 => "0000000000000000",
28251 => "0000000000000000",28252 => "0000000000000000",
28253 => "0000000000000000",28254 => "0000000000000000",
28255 => "0000000000000000",28256 => "0000000000000000",
28257 => "0000000000000000",28258 => "0000000000000000",
28259 => "0000000000000000",28260 => "0000000000000000",
28261 => "0000000000000000",28262 => "0000000000000000",
28263 => "0000000000000000",28264 => "0000000000000000",
28265 => "0000000000000000",28266 => "0000000000000000",
28267 => "0000000000000000",28268 => "0000000000000000",
28269 => "0000000000000000",28270 => "0000000000000000",
28271 => "0000000000000000",28272 => "0000000000000000",
28273 => "0000000000000000",28274 => "0000000000000000",
28275 => "0000000000000000",28276 => "0000000000000000",
28277 => "0000000000000000",28278 => "0000000000000000",
28279 => "0000000000000000",28280 => "0000000000000000",
28281 => "0000000000000000",28282 => "0000000000000000",
28283 => "0000000000000000",28284 => "0000000000000000",
28285 => "0000000000000000",28286 => "0000000000000000",
28287 => "0000000000000000",28288 => "0000000000000000",
28289 => "0000000000000000",28290 => "0000000000000000",
28291 => "0000000000000000",28292 => "0000000000000000",
28293 => "0000000000000000",28294 => "0000000000000000",
28295 => "0000000000000000",28296 => "0000000000000000",
28297 => "0000000000000000",28298 => "0000000000000000",
28299 => "0000000000000000",28300 => "0000000000000000",
28301 => "0000000000000000",28302 => "0000000000000000",
28303 => "0000000000000000",28304 => "0000000000000000",
28305 => "0000000000000000",28306 => "0000000000000000",
28307 => "0000000000000000",28308 => "0000000000000000",
28309 => "0000000000000000",28310 => "0000000000000000",
28311 => "0000000000000000",28312 => "0000000000000000",
28313 => "0000000000000000",28314 => "0000000000000000",
28315 => "0000000000000000",28316 => "0000000000000000",
28317 => "0000000000000000",28318 => "0000000000000000",
28319 => "0000000000000000",28320 => "0000000000000000",
28321 => "0000000000000000",28322 => "0000000000000000",
28323 => "0000000000000000",28324 => "0000000000000000",
28325 => "0000000000000000",28326 => "0000000000000000",
28327 => "0000000000000000",28328 => "0000000000000000",
28329 => "0000000000000000",28330 => "0000000000000000",
28331 => "0000000000000000",28332 => "0000000000000000",
28333 => "0000000000000000",28334 => "0000000000000000",
28335 => "0000000000000000",28336 => "0000000000000000",
28337 => "0000000000000000",28338 => "0000000000000000",
28339 => "0000000000000000",28340 => "0000000000000000",
28341 => "0000000000000000",28342 => "0000000000000000",
28343 => "0000000000000000",28344 => "0000000000000000",
28345 => "0000000000000000",28346 => "0000000000000000",
28347 => "0000000000000000",28348 => "0000000000000000",
28349 => "0000000000000000",28350 => "0000000000000000",
28351 => "0000000000000000",28352 => "0000000000000000",
28353 => "0000000000000000",28354 => "0000000000000000",
28355 => "0000000000000000",28356 => "0000000000000000",
28357 => "0000000000000000",28358 => "0000000000000000",
28359 => "0000000000000000",28360 => "0000000000000000",
28361 => "0000000000000000",28362 => "0000000000000000",
28363 => "0000000000000000",28364 => "0000000000000000",
28365 => "0000000000000000",28366 => "0000000000000000",
28367 => "0000000000000000",28368 => "0000000000000000",
28369 => "0000000000000000",28370 => "0000000000000000",
28371 => "0000000000000000",28372 => "0000000000000000",
28373 => "0000000000000000",28374 => "0000000000000000",
28375 => "0000000000000000",28376 => "0000000000000000",
28377 => "0000000000000000",28378 => "0000000000000000",
28379 => "0000000000000000",28380 => "0000000000000000",
28381 => "0000000000000000",28382 => "0000000000000000",
28383 => "0000000000000000",28384 => "0000000000000000",
28385 => "0000000000000000",28386 => "0000000000000000",
28387 => "0000000000000000",28388 => "0000000000000000",
28389 => "0000000000000000",28390 => "0000000000000000",
28391 => "0000000000000000",28392 => "0000000000000000",
28393 => "0000000000000000",28394 => "0000000000000000",
28395 => "0000000000000000",28396 => "0000000000000000",
28397 => "0000000000000000",28398 => "0000000000000000",
28399 => "0000000000000000",28400 => "0000000000000000",
28401 => "0000000000000000",28402 => "0000000000000000",
28403 => "0000000000000000",28404 => "0000000000000000",
28405 => "0000000000000000",28406 => "0000000000000000",
28407 => "0000000000000000",28408 => "0000000000000000",
28409 => "0000000000000000",28410 => "0000000000000000",
28411 => "0000000000000000",28412 => "0000000000000000",
28413 => "0000000000000000",28414 => "0000000000000000",
28415 => "0000000000000000",28416 => "0000000000000000",
28417 => "0000000000000000",28418 => "0000000000000000",
28419 => "0000000000000000",28420 => "0000000000000000",
28421 => "0000000000000000",28422 => "0000000000000000",
28423 => "0000000000000000",28424 => "0000000000000000",
28425 => "0000000000000000",28426 => "0000000000000000",
28427 => "0000000000000000",28428 => "0000000000000000",
28429 => "0000000000000000",28430 => "0000000000000000",
28431 => "0000000000000000",28432 => "0000000000000000",
28433 => "0000000000000000",28434 => "0000000000000000",
28435 => "0000000000000000",28436 => "0000000000000000",
28437 => "0000000000000000",28438 => "0000000000000000",
28439 => "0000000000000000",28440 => "0000000000000000",
28441 => "0000000000000000",28442 => "0000000000000000",
28443 => "0000000000000000",28444 => "0000000000000000",
28445 => "0000000000000000",28446 => "0000000000000000",
28447 => "0000000000000000",28448 => "0000000000000000",
28449 => "0000000000000000",28450 => "0000000000000000",
28451 => "0000000000000000",28452 => "0000000000000000",
28453 => "0000000000000000",28454 => "0000000000000000",
28455 => "0000000000000000",28456 => "0000000000000000",
28457 => "0000000000000000",28458 => "0000000000000000",
28459 => "0000000000000000",28460 => "0000000000000000",
28461 => "0000000000000000",28462 => "0000000000000000",
28463 => "0000000000000000",28464 => "0000000000000000",
28465 => "0000000000000000",28466 => "0000000000000000",
28467 => "0000000000000000",28468 => "0000000000000000",
28469 => "0000000000000000",28470 => "0000000000000000",
28471 => "0000000000000000",28472 => "0000000000000000",
28473 => "0000000000000000",28474 => "0000000000000000",
28475 => "0000000000000000",28476 => "0000000000000000",
28477 => "0000000000000000",28478 => "0000000000000000",
28479 => "0000000000000000",28480 => "0000000000000000",
28481 => "0000000000000000",28482 => "0000000000000000",
28483 => "0000000000000000",28484 => "0000000000000000",
28485 => "0000000000000000",28486 => "0000000000000000",
28487 => "0000000000000000",28488 => "0000000000000000",
28489 => "0000000000000000",28490 => "0000000000000000",
28491 => "0000000000000000",28492 => "0000000000000000",
28493 => "0000000000000000",28494 => "0000000000000000",
28495 => "0000000000000000",28496 => "0000000000000000",
28497 => "0000000000000000",28498 => "0000000000000000",
28499 => "0000000000000000",28500 => "0000000000000000",
28501 => "0000000000000000",28502 => "0000000000000000",
28503 => "0000000000000000",28504 => "0000000000000000",
28505 => "0000000000000000",28506 => "0000000000000000",
28507 => "0000000000000000",28508 => "0000000000000000",
28509 => "0000000000000000",28510 => "0000000000000000",
28511 => "0000000000000000",28512 => "0000000000000000",
28513 => "0000000000000000",28514 => "0000000000000000",
28515 => "0000000000000000",28516 => "0000000000000000",
28517 => "0000000000000000",28518 => "0000000000000000",
28519 => "0000000000000000",28520 => "0000000000000000",
28521 => "0000000000000000",28522 => "0000000000000000",
28523 => "0000000000000000",28524 => "0000000000000000",
28525 => "0000000000000000",28526 => "0000000000000000",
28527 => "0000000000000000",28528 => "0000000000000000",
28529 => "0000000000000000",28530 => "0000000000000000",
28531 => "0000000000000000",28532 => "0000000000000000",
28533 => "0000000000000000",28534 => "0000000000000000",
28535 => "0000000000000000",28536 => "0000000000000000",
28537 => "0000000000000000",28538 => "0000000000000000",
28539 => "0000000000000000",28540 => "0000000000000000",
28541 => "0000000000000000",28542 => "0000000000000000",
28543 => "0000000000000000",28544 => "0000000000000000",
28545 => "0000000000000000",28546 => "0000000000000000",
28547 => "0000000000000000",28548 => "0000000000000000",
28549 => "0000000000000000",28550 => "0000000000000000",
28551 => "0000000000000000",28552 => "0000000000000000",
28553 => "0000000000000000",28554 => "0000000000000000",
28555 => "0000000000000000",28556 => "0000000000000000",
28557 => "0000000000000000",28558 => "0000000000000000",
28559 => "0000000000000000",28560 => "0000000000000000",
28561 => "0000000000000000",28562 => "0000000000000000",
28563 => "0000000000000000",28564 => "0000000000000000",
28565 => "0000000000000000",28566 => "0000000000000000",
28567 => "0000000000000000",28568 => "0000000000000000",
28569 => "0000000000000000",28570 => "0000000000000000",
28571 => "0000000000000000",28572 => "0000000000000000",
28573 => "0000000000000000",28574 => "0000000000000000",
28575 => "0000000000000000",28576 => "0000000000000000",
28577 => "0000000000000000",28578 => "0000000000000000",
28579 => "0000000000000000",28580 => "0000000000000000",
28581 => "0000000000000000",28582 => "0000000000000000",
28583 => "0000000000000000",28584 => "0000000000000000",
28585 => "0000000000000000",28586 => "0000000000000000",
28587 => "0000000000000000",28588 => "0000000000000000",
28589 => "0000000000000000",28590 => "0000000000000000",
28591 => "0000000000000000",28592 => "0000000000000000",
28593 => "0000000000000000",28594 => "0000000000000000",
28595 => "0000000000000000",28596 => "0000000000000000",
28597 => "0000000000000000",28598 => "0000000000000000",
28599 => "0000000000000000",28600 => "0000000000000000",
28601 => "0000000000000000",28602 => "0000000000000000",
28603 => "0000000000000000",28604 => "0000000000000000",
28605 => "0000000000000000",28606 => "0000000000000000",
28607 => "0000000000000000",28608 => "0000000000000000",
28609 => "0000000000000000",28610 => "0000000000000000",
28611 => "0000000000000000",28612 => "0000000000000000",
28613 => "0000000000000000",28614 => "0000000000000000",
28615 => "0000000000000000",28616 => "0000000000000000",
28617 => "0000000000000000",28618 => "0000000000000000",
28619 => "0000000000000000",28620 => "0000000000000000",
28621 => "0000000000000000",28622 => "0000000000000000",
28623 => "0000000000000000",28624 => "0000000000000000",
28625 => "0000000000000000",28626 => "0000000000000000",
28627 => "0000000000000000",28628 => "0000000000000000",
28629 => "0000000000000000",28630 => "0000000000000000",
28631 => "0000000000000000",28632 => "0000000000000000",
28633 => "0000000000000000",28634 => "0000000000000000",
28635 => "0000000000000000",28636 => "0000000000000000",
28637 => "0000000000000000",28638 => "0000000000000000",
28639 => "0000000000000000",28640 => "0000000000000000",
28641 => "0000000000000000",28642 => "0000000000000000",
28643 => "0000000000000000",28644 => "0000000000000000",
28645 => "0000000000000000",28646 => "0000000000000000",
28647 => "0000000000000000",28648 => "0000000000000000",
28649 => "0000000000000000",28650 => "0000000000000000",
28651 => "0000000000000000",28652 => "0000000000000000",
28653 => "0000000000000000",28654 => "0000000000000000",
28655 => "0000000000000000",28656 => "0000000000000000",
28657 => "0000000000000000",28658 => "0000000000000000",
28659 => "0000000000000000",28660 => "0000000000000000",
28661 => "0000000000000000",28662 => "0000000000000000",
28663 => "0000000000000000",28664 => "0000000000000000",
28665 => "0000000000000000",28666 => "0000000000000000",
28667 => "0000000000000000",28668 => "0000000000000000",
28669 => "0000000000000000",28670 => "0000000000000000",
28671 => "0000000000000000",28672 => "0000000000000000",
28673 => "0000000000000000",28674 => "0000000000000000",
28675 => "0000000000000000",28676 => "0000000000000000",
28677 => "0000000000000000",28678 => "0000000000000000",
28679 => "0000000000000000",28680 => "0000000000000000",
28681 => "0000000000000000",28682 => "0000000000000000",
28683 => "0000000000000000",28684 => "0000000000000000",
28685 => "0000000000000000",28686 => "0000000000000000",
28687 => "0000000000000000",28688 => "0000000000000000",
28689 => "0000000000000000",28690 => "0000000000000000",
28691 => "0000000000000000",28692 => "0000000000000000",
28693 => "0000000000000000",28694 => "0000000000000000",
28695 => "0000000000000000",28696 => "0000000000000000",
28697 => "0000000000000000",28698 => "0000000000000000",
28699 => "0000000000000000",28700 => "0000000000000000",
28701 => "0000000000000000",28702 => "0000000000000000",
28703 => "0000000000000000",28704 => "0000000000000000",
28705 => "0000000000000000",28706 => "0000000000000000",
28707 => "0000000000000000",28708 => "0000000000000000",
28709 => "0000000000000000",28710 => "0000000000000000",
28711 => "0000000000000000",28712 => "0000000000000000",
28713 => "0000000000000000",28714 => "0000000000000000",
28715 => "0000000000000000",28716 => "0000000000000000",
28717 => "0000000000000000",28718 => "0000000000000000",
28719 => "0000000000000000",28720 => "0000000000000000",
28721 => "0000000000000000",28722 => "0000000000000000",
28723 => "0000000000000000",28724 => "0000000000000000",
28725 => "0000000000000000",28726 => "0000000000000000",
28727 => "0000000000000000",28728 => "0000000000000000",
28729 => "0000000000000000",28730 => "0000000000000000",
28731 => "0000000000000000",28732 => "0000000000000000",
28733 => "0000000000000000",28734 => "0000000000000000",
28735 => "0000000000000000",28736 => "0000000000000000",
28737 => "0000000000000000",28738 => "0000000000000000",
28739 => "0000000000000000",28740 => "0000000000000000",
28741 => "0000000000000000",28742 => "0000000000000000",
28743 => "0000000000000000",28744 => "0000000000000000",
28745 => "0000000000000000",28746 => "0000000000000000",
28747 => "0000000000000000",28748 => "0000000000000000",
28749 => "0000000000000000",28750 => "0000000000000000",
28751 => "0000000000000000",28752 => "0000000000000000",
28753 => "0000000000000000",28754 => "0000000000000000",
28755 => "0000000000000000",28756 => "0000000000000000",
28757 => "0000000000000000",28758 => "0000000000000000",
28759 => "0000000000000000",28760 => "0000000000000000",
28761 => "0000000000000000",28762 => "0000000000000000",
28763 => "0000000000000000",28764 => "0000000000000000",
28765 => "0000000000000000",28766 => "0000000000000000",
28767 => "0000000000000000",28768 => "0000000000000000",
28769 => "0000000000000000",28770 => "0000000000000000",
28771 => "0000000000000000",28772 => "0000000000000000",
28773 => "0000000000000000",28774 => "0000000000000000",
28775 => "0000000000000000",28776 => "0000000000000000",
28777 => "0000000000000000",28778 => "0000000000000000",
28779 => "0000000000000000",28780 => "0000000000000000",
28781 => "0000000000000000",28782 => "0000000000000000",
28783 => "0000000000000000",28784 => "0000000000000000",
28785 => "0000000000000000",28786 => "0000000000000000",
28787 => "0000000000000000",28788 => "0000000000000000",
28789 => "0000000000000000",28790 => "0000000000000000",
28791 => "0000000000000000",28792 => "0000000000000000",
28793 => "0000000000000000",28794 => "0000000000000000",
28795 => "0000000000000000",28796 => "0000000000000000",
28797 => "0000000000000000",28798 => "0000000000000000",
28799 => "0000000000000000",28800 => "0000000000000000",
28801 => "0000000000000000",28802 => "0000000000000000",
28803 => "0000000000000000",28804 => "0000000000000000",
28805 => "0000000000000000",28806 => "0000000000000000",
28807 => "0000000000000000",28808 => "0000000000000000",
28809 => "0000000000000000",28810 => "0000000000000000",
28811 => "0000000000000000",28812 => "0000000000000000",
28813 => "0000000000000000",28814 => "0000000000000000",
28815 => "0000000000000000",28816 => "0000000000000000",
28817 => "0000000000000000",28818 => "0000000000000000",
28819 => "0000000000000000",28820 => "0000000000000000",
28821 => "0000000000000000",28822 => "0000000000000000",
28823 => "0000000000000000",28824 => "0000000000000000",
28825 => "0000000000000000",28826 => "0000000000000000",
28827 => "0000000000000000",28828 => "0000000000000000",
28829 => "0000000000000000",28830 => "0000000000000000",
28831 => "0000000000000000",28832 => "0000000000000000",
28833 => "0000000000000000",28834 => "0000000000000000",
28835 => "0000000000000000",28836 => "0000000000000000",
28837 => "0000000000000000",28838 => "0000000000000000",
28839 => "0000000000000000",28840 => "0000000000000000",
28841 => "0000000000000000",28842 => "0000000000000000",
28843 => "0000000000000000",28844 => "0000000000000000",
28845 => "0000000000000000",28846 => "0000000000000000",
28847 => "0000000000000000",28848 => "0000000000000000",
28849 => "0000000000000000",28850 => "0000000000000000",
28851 => "0000000000000000",28852 => "0000000000000000",
28853 => "0000000000000000",28854 => "0000000000000000",
28855 => "0000000000000000",28856 => "0000000000000000",
28857 => "0000000000000000",28858 => "0000000000000000",
28859 => "0000000000000000",28860 => "0000000000000000",
28861 => "0000000000000000",28862 => "0000000000000000",
28863 => "0000000000000000",28864 => "0000000000000000",
28865 => "0000000000000000",28866 => "0000000000000000",
28867 => "0000000000000000",28868 => "0000000000000000",
28869 => "0000000000000000",28870 => "0000000000000000",
28871 => "0000000000000000",28872 => "0000000000000000",
28873 => "0000000000000000",28874 => "0000000000000000",
28875 => "0000000000000000",28876 => "0000000000000000",
28877 => "0000000000000000",28878 => "0000000000000000",
28879 => "0000000000000000",28880 => "0000000000000000",
28881 => "0000000000000000",28882 => "0000000000000000",
28883 => "0000000000000000",28884 => "0000000000000000",
28885 => "0000000000000000",28886 => "0000000000000000",
28887 => "0000000000000000",28888 => "0000000000000000",
28889 => "0000000000000000",28890 => "0000000000000000",
28891 => "0000000000000000",28892 => "0000000000000000",
28893 => "0000000000000000",28894 => "0000000000000000",
28895 => "0000000000000000",28896 => "0000000000000000",
28897 => "0000000000000000",28898 => "0000000000000000",
28899 => "0000000000000000",28900 => "0000000000000000",
28901 => "0000000000000000",28902 => "0000000000000000",
28903 => "0000000000000000",28904 => "0000000000000000",
28905 => "0000000000000000",28906 => "0000000000000000",
28907 => "0000000000000000",28908 => "0000000000000000",
28909 => "0000000000000000",28910 => "0000000000000000",
28911 => "0000000000000000",28912 => "0000000000000000",
28913 => "0000000000000000",28914 => "0000000000000000",
28915 => "0000000000000000",28916 => "0000000000000000",
28917 => "0000000000000000",28918 => "0000000000000000",
28919 => "0000000000000000",28920 => "0000000000000000",
28921 => "0000000000000000",28922 => "0000000000000000",
28923 => "0000000000000000",28924 => "0000000000000000",
28925 => "0000000000000000",28926 => "0000000000000000",
28927 => "0000000000000000",28928 => "0000000000000000",
28929 => "0000000000000000",28930 => "0000000000000000",
28931 => "0000000000000000",28932 => "0000000000000000",
28933 => "0000000000000000",28934 => "0000000000000000",
28935 => "0000000000000000",28936 => "0000000000000000",
28937 => "0000000000000000",28938 => "0000000000000000",
28939 => "0000000000000000",28940 => "0000000000000000",
28941 => "0000000000000000",28942 => "0000000000000000",
28943 => "0000000000000000",28944 => "0000000000000000",
28945 => "0000000000000000",28946 => "0000000000000000",
28947 => "0000000000000000",28948 => "0000000000000000",
28949 => "0000000000000000",28950 => "0000000000000000",
28951 => "0000000000000000",28952 => "0000000000000000",
28953 => "0000000000000000",28954 => "0000000000000000",
28955 => "0000000000000000",28956 => "0000000000000000",
28957 => "0000000000000000",28958 => "0000000000000000",
28959 => "0000000000000000",28960 => "0000000000000000",
28961 => "0000000000000000",28962 => "0000000000000000",
28963 => "0000000000000000",28964 => "0000000000000000",
28965 => "0000000000000000",28966 => "0000000000000000",
28967 => "0000000000000000",28968 => "0000000000000000",
28969 => "0000000000000000",28970 => "0000000000000000",
28971 => "0000000000000000",28972 => "0000000000000000",
28973 => "0000000000000000",28974 => "0000000000000000",
28975 => "0000000000000000",28976 => "0000000000000000",
28977 => "0000000000000000",28978 => "0000000000000000",
28979 => "0000000000000000",28980 => "0000000000000000",
28981 => "0000000000000000",28982 => "0000000000000000",
28983 => "0000000000000000",28984 => "0000000000000000",
28985 => "0000000000000000",28986 => "0000000000000000",
28987 => "0000000000000000",28988 => "0000000000000000",
28989 => "0000000000000000",28990 => "0000000000000000",
28991 => "0000000000000000",28992 => "0000000000000000",
28993 => "0000000000000000",28994 => "0000000000000000",
28995 => "0000000000000000",28996 => "0000000000000000",
28997 => "0000000000000000",28998 => "0000000000000000",
28999 => "0000000000000000",29000 => "0000000000000000",
29001 => "0000000000000000",29002 => "0000000000000000",
29003 => "0000000000000000",29004 => "0000000000000000",
29005 => "0000000000000000",29006 => "0000000000000000",
29007 => "0000000000000000",29008 => "0000000000000000",
29009 => "0000000000000000",29010 => "0000000000000000",
29011 => "0000000000000000",29012 => "0000000000000000",
29013 => "0000000000000000",29014 => "0000000000000000",
29015 => "0000000000000000",29016 => "0000000000000000",
29017 => "0000000000000000",29018 => "0000000000000000",
29019 => "0000000000000000",29020 => "0000000000000000",
29021 => "0000000000000000",29022 => "0000000000000000",
29023 => "0000000000000000",29024 => "0000000000000000",
29025 => "0000000000000000",29026 => "0000000000000000",
29027 => "0000000000000000",29028 => "0000000000000000",
29029 => "0000000000000000",29030 => "0000000000000000",
29031 => "0000000000000000",29032 => "0000000000000000",
29033 => "0000000000000000",29034 => "0000000000000000",
29035 => "0000000000000000",29036 => "0000000000000000",
29037 => "0000000000000000",29038 => "0000000000000000",
29039 => "0000000000000000",29040 => "0000000000000000",
29041 => "0000000000000000",29042 => "0000000000000000",
29043 => "0000000000000000",29044 => "0000000000000000",
29045 => "0000000000000000",29046 => "0000000000000000",
29047 => "0000000000000000",29048 => "0000000000000000",
29049 => "0000000000000000",29050 => "0000000000000000",
29051 => "0000000000000000",29052 => "0000000000000000",
29053 => "0000000000000000",29054 => "0000000000000000",
29055 => "0000000000000000",29056 => "0000000000000000",
29057 => "0000000000000000",29058 => "0000000000000000",
29059 => "0000000000000000",29060 => "0000000000000000",
29061 => "0000000000000000",29062 => "0000000000000000",
29063 => "0000000000000000",29064 => "0000000000000000",
29065 => "0000000000000000",29066 => "0000000000000000",
29067 => "0000000000000000",29068 => "0000000000000000",
29069 => "0000000000000000",29070 => "0000000000000000",
29071 => "0000000000000000",29072 => "0000000000000000",
29073 => "0000000000000000",29074 => "0000000000000000",
29075 => "0000000000000000",29076 => "0000000000000000",
29077 => "0000000000000000",29078 => "0000000000000000",
29079 => "0000000000000000",29080 => "0000000000000000",
29081 => "0000000000000000",29082 => "0000000000000000",
29083 => "0000000000000000",29084 => "0000000000000000",
29085 => "0000000000000000",29086 => "0000000000000000",
29087 => "0000000000000000",29088 => "0000000000000000",
29089 => "0000000000000000",29090 => "0000000000000000",
29091 => "0000000000000000",29092 => "0000000000000000",
29093 => "0000000000000000",29094 => "0000000000000000",
29095 => "0000000000000000",29096 => "0000000000000000",
29097 => "0000000000000000",29098 => "0000000000000000",
29099 => "0000000000000000",29100 => "0000000000000000",
29101 => "0000000000000000",29102 => "0000000000000000",
29103 => "0000000000000000",29104 => "0000000000000000",
29105 => "0000000000000000",29106 => "0000000000000000",
29107 => "0000000000000000",29108 => "0000000000000000",
29109 => "0000000000000000",29110 => "0000000000000000",
29111 => "0000000000000000",29112 => "0000000000000000",
29113 => "0000000000000000",29114 => "0000000000000000",
29115 => "0000000000000000",29116 => "0000000000000000",
29117 => "0000000000000000",29118 => "0000000000000000",
29119 => "0000000000000000",29120 => "0000000000000000",
29121 => "0000000000000000",29122 => "0000000000000000",
29123 => "0000000000000000",29124 => "0000000000000000",
29125 => "0000000000000000",29126 => "0000000000000000",
29127 => "0000000000000000",29128 => "0000000000000000",
29129 => "0000000000000000",29130 => "0000000000000000",
29131 => "0000000000000000",29132 => "0000000000000000",
29133 => "0000000000000000",29134 => "0000000000000000",
29135 => "0000000000000000",29136 => "0000000000000000",
29137 => "0000000000000000",29138 => "0000000000000000",
29139 => "0000000000000000",29140 => "0000000000000000",
29141 => "0000000000000000",29142 => "0000000000000000",
29143 => "0000000000000000",29144 => "0000000000000000",
29145 => "0000000000000000",29146 => "0000000000000000",
29147 => "0000000000000000",29148 => "0000000000000000",
29149 => "0000000000000000",29150 => "0000000000000000",
29151 => "0000000000000000",29152 => "0000000000000000",
29153 => "0000000000000000",29154 => "0000000000000000",
29155 => "0000000000000000",29156 => "0000000000000000",
29157 => "0000000000000000",29158 => "0000000000000000",
29159 => "0000000000000000",29160 => "0000000000000000",
29161 => "0000000000000000",29162 => "0000000000000000",
29163 => "0000000000000000",29164 => "0000000000000000",
29165 => "0000000000000000",29166 => "0000000000000000",
29167 => "0000000000000000",29168 => "0000000000000000",
29169 => "0000000000000000",29170 => "0000000000000000",
29171 => "0000000000000000",29172 => "0000000000000000",
29173 => "0000000000000000",29174 => "0000000000000000",
29175 => "0000000000000000",29176 => "0000000000000000",
29177 => "0000000000000000",29178 => "0000000000000000",
29179 => "0000000000000000",29180 => "0000000000000000",
29181 => "0000000000000000",29182 => "0000000000000000",
29183 => "0000000000000000",29184 => "0000000000000000",
29185 => "0000000000000000",29186 => "0000000000000000",
29187 => "0000000000000000",29188 => "0000000000000000",
29189 => "0000000000000000",29190 => "0000000000000000",
29191 => "0000000000000000",29192 => "0000000000000000",
29193 => "0000000000000000",29194 => "0000000000000000",
29195 => "0000000000000000",29196 => "0000000000000000",
29197 => "0000000000000000",29198 => "0000000000000000",
29199 => "0000000000000000",29200 => "0000000000000000",
29201 => "0000000000000000",29202 => "0000000000000000",
29203 => "0000000000000000",29204 => "0000000000000000",
29205 => "0000000000000000",29206 => "0000000000000000",
29207 => "0000000000000000",29208 => "0000000000000000",
29209 => "0000000000000000",29210 => "0000000000000000",
29211 => "0000000000000000",29212 => "0000000000000000",
29213 => "0000000000000000",29214 => "0000000000000000",
29215 => "0000000000000000",29216 => "0000000000000000",
29217 => "0000000000000000",29218 => "0000000000000000",
29219 => "0000000000000000",29220 => "0000000000000000",
29221 => "0000000000000000",29222 => "0000000000000000",
29223 => "0000000000000000",29224 => "0000000000000000",
29225 => "0000000000000000",29226 => "0000000000000000",
29227 => "0000000000000000",29228 => "0000000000000000",
29229 => "0000000000000000",29230 => "0000000000000000",
29231 => "0000000000000000",29232 => "0000000000000000",
29233 => "0000000000000000",29234 => "0000000000000000",
29235 => "0000000000000000",29236 => "0000000000000000",
29237 => "0000000000000000",29238 => "0000000000000000",
29239 => "0000000000000000",29240 => "0000000000000000",
29241 => "0000000000000000",29242 => "0000000000000000",
29243 => "0000000000000000",29244 => "0000000000000000",
29245 => "0000000000000000",29246 => "0000000000000000",
29247 => "0000000000000000",29248 => "0000000000000000",
29249 => "0000000000000000",29250 => "0000000000000000",
29251 => "0000000000000000",29252 => "0000000000000000",
29253 => "0000000000000000",29254 => "0000000000000000",
29255 => "0000000000000000",29256 => "0000000000000000",
29257 => "0000000000000000",29258 => "0000000000000000",
29259 => "0000000000000000",29260 => "0000000000000000",
29261 => "0000000000000000",29262 => "0000000000000000",
29263 => "0000000000000000",29264 => "0000000000000000",
29265 => "0000000000000000",29266 => "0000000000000000",
29267 => "0000000000000000",29268 => "0000000000000000",
29269 => "0000000000000000",29270 => "0000000000000000",
29271 => "0000000000000000",29272 => "0000000000000000",
29273 => "0000000000000000",29274 => "0000000000000000",
29275 => "0000000000000000",29276 => "0000000000000000",
29277 => "0000000000000000",29278 => "0000000000000000",
29279 => "0000000000000000",29280 => "0000000000000000",
29281 => "0000000000000000",29282 => "0000000000000000",
29283 => "0000000000000000",29284 => "0000000000000000",
29285 => "0000000000000000",29286 => "0000000000000000",
29287 => "0000000000000000",29288 => "0000000000000000",
29289 => "0000000000000000",29290 => "0000000000000000",
29291 => "0000000000000000",29292 => "0000000000000000",
29293 => "0000000000000000",29294 => "0000000000000000",
29295 => "0000000000000000",29296 => "0000000000000000",
29297 => "0000000000000000",29298 => "0000000000000000",
29299 => "0000000000000000",29300 => "0000000000000000",
29301 => "0000000000000000",29302 => "0000000000000000",
29303 => "0000000000000000",29304 => "0000000000000000",
29305 => "0000000000000000",29306 => "0000000000000000",
29307 => "0000000000000000",29308 => "0000000000000000",
29309 => "0000000000000000",29310 => "0000000000000000",
29311 => "0000000000000000",29312 => "0000000000000000",
29313 => "0000000000000000",29314 => "0000000000000000",
29315 => "0000000000000000",29316 => "0000000000000000",
29317 => "0000000000000000",29318 => "0000000000000000",
29319 => "0000000000000000",29320 => "0000000000000000",
29321 => "0000000000000000",29322 => "0000000000000000",
29323 => "0000000000000000",29324 => "0000000000000000",
29325 => "0000000000000000",29326 => "0000000000000000",
29327 => "0000000000000000",29328 => "0000000000000000",
29329 => "0000000000000000",29330 => "0000000000000000",
29331 => "0000000000000000",29332 => "0000000000000000",
29333 => "0000000000000000",29334 => "0000000000000000",
29335 => "0000000000000000",29336 => "0000000000000000",
29337 => "0000000000000000",29338 => "0000000000000000",
29339 => "0000000000000000",29340 => "0000000000000000",
29341 => "0000000000000000",29342 => "0000000000000000",
29343 => "0000000000000000",29344 => "0000000000000000",
29345 => "0000000000000000",29346 => "0000000000000000",
29347 => "0000000000000000",29348 => "0000000000000000",
29349 => "0000000000000000",29350 => "0000000000000000",
29351 => "0000000000000000",29352 => "0000000000000000",
29353 => "0000000000000000",29354 => "0000000000000000",
29355 => "0000000000000000",29356 => "0000000000000000",
29357 => "0000000000000000",29358 => "0000000000000000",
29359 => "0000000000000000",29360 => "0000000000000000",
29361 => "0000000000000000",29362 => "0000000000000000",
29363 => "0000000000000000",29364 => "0000000000000000",
29365 => "0000000000000000",29366 => "0000000000000000",
29367 => "0000000000000000",29368 => "0000000000000000",
29369 => "0000000000000000",29370 => "0000000000000000",
29371 => "0000000000000000",29372 => "0000000000000000",
29373 => "0000000000000000",29374 => "0000000000000000",
29375 => "0000000000000000",29376 => "0000000000000000",
29377 => "0000000000000000",29378 => "0000000000000000",
29379 => "0000000000000000",29380 => "0000000000000000",
29381 => "0000000000000000",29382 => "0000000000000000",
29383 => "0000000000000000",29384 => "0000000000000000",
29385 => "0000000000000000",29386 => "0000000000000000",
29387 => "0000000000000000",29388 => "0000000000000000",
29389 => "0000000000000000",29390 => "0000000000000000",
29391 => "0000000000000000",29392 => "0000000000000000",
29393 => "0000000000000000",29394 => "0000000000000000",
29395 => "0000000000000000",29396 => "0000000000000000",
29397 => "0000000000000000",29398 => "0000000000000000",
29399 => "0000000000000000",29400 => "0000000000000000",
29401 => "0000000000000000",29402 => "0000000000000000",
29403 => "0000000000000000",29404 => "0000000000000000",
29405 => "0000000000000000",29406 => "0000000000000000",
29407 => "0000000000000000",29408 => "0000000000000000",
29409 => "0000000000000000",29410 => "0000000000000000",
29411 => "0000000000000000",29412 => "0000000000000000",
29413 => "0000000000000000",29414 => "0000000000000000",
29415 => "0000000000000000",29416 => "0000000000000000",
29417 => "0000000000000000",29418 => "0000000000000000",
29419 => "0000000000000000",29420 => "0000000000000000",
29421 => "0000000000000000",29422 => "0000000000000000",
29423 => "0000000000000000",29424 => "0000000000000000",
29425 => "0000000000000000",29426 => "0000000000000000",
29427 => "0000000000000000",29428 => "0000000000000000",
29429 => "0000000000000000",29430 => "0000000000000000",
29431 => "0000000000000000",29432 => "0000000000000000",
29433 => "0000000000000000",29434 => "0000000000000000",
29435 => "0000000000000000",29436 => "0000000000000000",
29437 => "0000000000000000",29438 => "0000000000000000",
29439 => "0000000000000000",29440 => "0000000000000000",
29441 => "0000000000000000",29442 => "0000000000000000",
29443 => "0000000000000000",29444 => "0000000000000000",
29445 => "0000000000000000",29446 => "0000000000000000",
29447 => "0000000000000000",29448 => "0000000000000000",
29449 => "0000000000000000",29450 => "0000000000000000",
29451 => "0000000000000000",29452 => "0000000000000000",
29453 => "0000000000000000",29454 => "0000000000000000",
29455 => "0000000000000000",29456 => "0000000000000000",
29457 => "0000000000000000",29458 => "0000000000000000",
29459 => "0000000000000000",29460 => "0000000000000000",
29461 => "0000000000000000",29462 => "0000000000000000",
29463 => "0000000000000000",29464 => "0000000000000000",
29465 => "0000000000000000",29466 => "0000000000000000",
29467 => "0000000000000000",29468 => "0000000000000000",
29469 => "0000000000000000",29470 => "0000000000000000",
29471 => "0000000000000000",29472 => "0000000000000000",
29473 => "0000000000000000",29474 => "0000000000000000",
29475 => "0000000000000000",29476 => "0000000000000000",
29477 => "0000000000000000",29478 => "0000000000000000",
29479 => "0000000000000000",29480 => "0000000000000000",
29481 => "0000000000000000",29482 => "0000000000000000",
29483 => "0000000000000000",29484 => "0000000000000000",
29485 => "0000000000000000",29486 => "0000000000000000",
29487 => "0000000000000000",29488 => "0000000000000000",
29489 => "0000000000000000",29490 => "0000000000000000",
29491 => "0000000000000000",29492 => "0000000000000000",
29493 => "0000000000000000",29494 => "0000000000000000",
29495 => "0000000000000000",29496 => "0000000000000000",
29497 => "0000000000000000",29498 => "0000000000000000",
29499 => "0000000000000000",29500 => "0000000000000000",
29501 => "0000000000000000",29502 => "0000000000000000",
29503 => "0000000000000000",29504 => "0000000000000000",
29505 => "0000000000000000",29506 => "0000000000000000",
29507 => "0000000000000000",29508 => "0000000000000000",
29509 => "0000000000000000",29510 => "0000000000000000",
29511 => "0000000000000000",29512 => "0000000000000000",
29513 => "0000000000000000",29514 => "0000000000000000",
29515 => "0000000000000000",29516 => "0000000000000000",
29517 => "0000000000000000",29518 => "0000000000000000",
29519 => "0000000000000000",29520 => "0000000000000000",
29521 => "0000000000000000",29522 => "0000000000000000",
29523 => "0000000000000000",29524 => "0000000000000000",
29525 => "0000000000000000",29526 => "0000000000000000",
29527 => "0000000000000000",29528 => "0000000000000000",
29529 => "0000000000000000",29530 => "0000000000000000",
29531 => "0000000000000000",29532 => "0000000000000000",
29533 => "0000000000000000",29534 => "0000000000000000",
29535 => "0000000000000000",29536 => "0000000000000000",
29537 => "0000000000000000",29538 => "0000000000000000",
29539 => "0000000000000000",29540 => "0000000000000000",
29541 => "0000000000000000",29542 => "0000000000000000",
29543 => "0000000000000000",29544 => "0000000000000000",
29545 => "0000000000000000",29546 => "0000000000000000",
29547 => "0000000000000000",29548 => "0000000000000000",
29549 => "0000000000000000",29550 => "0000000000000000",
29551 => "0000000000000000",29552 => "0000000000000000",
29553 => "0000000000000000",29554 => "0000000000000000",
29555 => "0000000000000000",29556 => "0000000000000000",
29557 => "0000000000000000",29558 => "0000000000000000",
29559 => "0000000000000000",29560 => "0000000000000000",
29561 => "0000000000000000",29562 => "0000000000000000",
29563 => "0000000000000000",29564 => "0000000000000000",
29565 => "0000000000000000",29566 => "0000000000000000",
29567 => "0000000000000000",29568 => "0000000000000000",
29569 => "0000000000000000",29570 => "0000000000000000",
29571 => "0000000000000000",29572 => "0000000000000000",
29573 => "0000000000000000",29574 => "0000000000000000",
29575 => "0000000000000000",29576 => "0000000000000000",
29577 => "0000000000000000",29578 => "0000000000000000",
29579 => "0000000000000000",29580 => "0000000000000000",
29581 => "0000000000000000",29582 => "0000000000000000",
29583 => "0000000000000000",29584 => "0000000000000000",
29585 => "0000000000000000",29586 => "0000000000000000",
29587 => "0000000000000000",29588 => "0000000000000000",
29589 => "0000000000000000",29590 => "0000000000000000",
29591 => "0000000000000000",29592 => "0000000000000000",
29593 => "0000000000000000",29594 => "0000000000000000",
29595 => "0000000000000000",29596 => "0000000000000000",
29597 => "0000000000000000",29598 => "0000000000000000",
29599 => "0000000000000000",29600 => "0000000000000000",
29601 => "0000000000000000",29602 => "0000000000000000",
29603 => "0000000000000000",29604 => "0000000000000000",
29605 => "0000000000000000",29606 => "0000000000000000",
29607 => "0000000000000000",29608 => "0000000000000000",
29609 => "0000000000000000",29610 => "0000000000000000",
29611 => "0000000000000000",29612 => "0000000000000000",
29613 => "0000000000000000",29614 => "0000000000000000",
29615 => "0000000000000000",29616 => "0000000000000000",
29617 => "0000000000000000",29618 => "0000000000000000",
29619 => "0000000000000000",29620 => "0000000000000000",
29621 => "0000000000000000",29622 => "0000000000000000",
29623 => "0000000000000000",29624 => "0000000000000000",
29625 => "0000000000000000",29626 => "0000000000000000",
29627 => "0000000000000000",29628 => "0000000000000000",
29629 => "0000000000000000",29630 => "0000000000000000",
29631 => "0000000000000000",29632 => "0000000000000000",
29633 => "0000000000000000",29634 => "0000000000000000",
29635 => "0000000000000000",29636 => "0000000000000000",
29637 => "0000000000000000",29638 => "0000000000000000",
29639 => "0000000000000000",29640 => "0000000000000000",
29641 => "0000000000000000",29642 => "0000000000000000",
29643 => "0000000000000000",29644 => "0000000000000000",
29645 => "0000000000000000",29646 => "0000000000000000",
29647 => "0000000000000000",29648 => "0000000000000000",
29649 => "0000000000000000",29650 => "0000000000000000",
29651 => "0000000000000000",29652 => "0000000000000000",
29653 => "0000000000000000",29654 => "0000000000000000",
29655 => "0000000000000000",29656 => "0000000000000000",
29657 => "0000000000000000",29658 => "0000000000000000",
29659 => "0000000000000000",29660 => "0000000000000000",
29661 => "0000000000000000",29662 => "0000000000000000",
29663 => "0000000000000000",29664 => "0000000000000000",
29665 => "0000000000000000",29666 => "0000000000000000",
29667 => "0000000000000000",29668 => "0000000000000000",
29669 => "0000000000000000",29670 => "0000000000000000",
29671 => "0000000000000000",29672 => "0000000000000000",
29673 => "0000000000000000",29674 => "0000000000000000",
29675 => "0000000000000000",29676 => "0000000000000000",
29677 => "0000000000000000",29678 => "0000000000000000",
29679 => "0000000000000000",29680 => "0000000000000000",
29681 => "0000000000000000",29682 => "0000000000000000",
29683 => "0000000000000000",29684 => "0000000000000000",
29685 => "0000000000000000",29686 => "0000000000000000",
29687 => "0000000000000000",29688 => "0000000000000000",
29689 => "0000000000000000",29690 => "0000000000000000",
29691 => "0000000000000000",29692 => "0000000000000000",
29693 => "0000000000000000",29694 => "0000000000000000",
29695 => "0000000000000000",29696 => "0000000000000000",
29697 => "0000000000000000",29698 => "0000000000000000",
29699 => "0000000000000000",29700 => "0000000000000000",
29701 => "0000000000000000",29702 => "0000000000000000",
29703 => "0000000000000000",29704 => "0000000000000000",
29705 => "0000000000000000",29706 => "0000000000000000",
29707 => "0000000000000000",29708 => "0000000000000000",
29709 => "0000000000000000",29710 => "0000000000000000",
29711 => "0000000000000000",29712 => "0000000000000000",
29713 => "0000000000000000",29714 => "0000000000000000",
29715 => "0000000000000000",29716 => "0000000000000000",
29717 => "0000000000000000",29718 => "0000000000000000",
29719 => "0000000000000000",29720 => "0000000000000000",
29721 => "0000000000000000",29722 => "0000000000000000",
29723 => "0000000000000000",29724 => "0000000000000000",
29725 => "0000000000000000",29726 => "0000000000000000",
29727 => "0000000000000000",29728 => "0000000000000000",
29729 => "0000000000000000",29730 => "0000000000000000",
29731 => "0000000000000000",29732 => "0000000000000000",
29733 => "0000000000000000",29734 => "0000000000000000",
29735 => "0000000000000000",29736 => "0000000000000000",
29737 => "0000000000000000",29738 => "0000000000000000",
29739 => "0000000000000000",29740 => "0000000000000000",
29741 => "0000000000000000",29742 => "0000000000000000",
29743 => "0000000000000000",29744 => "0000000000000000",
29745 => "0000000000000000",29746 => "0000000000000000",
29747 => "0000000000000000",29748 => "0000000000000000",
29749 => "0000000000000000",29750 => "0000000000000000",
29751 => "0000000000000000",29752 => "0000000000000000",
29753 => "0000000000000000",29754 => "0000000000000000",
29755 => "0000000000000000",29756 => "0000000000000000",
29757 => "0000000000000000",29758 => "0000000000000000",
29759 => "0000000000000000",29760 => "0000000000000000",
29761 => "0000000000000000",29762 => "0000000000000000",
29763 => "0000000000000000",29764 => "0000000000000000",
29765 => "0000000000000000",29766 => "0000000000000000",
29767 => "0000000000000000",29768 => "0000000000000000",
29769 => "0000000000000000",29770 => "0000000000000000",
29771 => "0000000000000000",29772 => "0000000000000000",
29773 => "0000000000000000",29774 => "0000000000000000",
29775 => "0000000000000000",29776 => "0000000000000000",
29777 => "0000000000000000",29778 => "0000000000000000",
29779 => "0000000000000000",29780 => "0000000000000000",
29781 => "0000000000000000",29782 => "0000000000000000",
29783 => "0000000000000000",29784 => "0000000000000000",
29785 => "0000000000000000",29786 => "0000000000000000",
29787 => "0000000000000000",29788 => "0000000000000000",
29789 => "0000000000000000",29790 => "0000000000000000",
29791 => "0000000000000000",29792 => "0000000000000000",
29793 => "0000000000000000",29794 => "0000000000000000",
29795 => "0000000000000000",29796 => "0000000000000000",
29797 => "0000000000000000",29798 => "0000000000000000",
29799 => "0000000000000000",29800 => "0000000000000000",
29801 => "0000000000000000",29802 => "0000000000000000",
29803 => "0000000000000000",29804 => "0000000000000000",
29805 => "0000000000000000",29806 => "0000000000000000",
29807 => "0000000000000000",29808 => "0000000000000000",
29809 => "0000000000000000",29810 => "0000000000000000",
29811 => "0000000000000000",29812 => "0000000000000000",
29813 => "0000000000000000",29814 => "0000000000000000",
29815 => "0000000000000000",29816 => "0000000000000000",
29817 => "0000000000000000",29818 => "0000000000000000",
29819 => "0000000000000000",29820 => "0000000000000000",
29821 => "0000000000000000",29822 => "0000000000000000",
29823 => "0000000000000000",29824 => "0000000000000000",
29825 => "0000000000000000",29826 => "0000000000000000",
29827 => "0000000000000000",29828 => "0000000000000000",
29829 => "0000000000000000",29830 => "0000000000000000",
29831 => "0000000000000000",29832 => "0000000000000000",
29833 => "0000000000000000",29834 => "0000000000000000",
29835 => "0000000000000000",29836 => "0000000000000000",
29837 => "0000000000000000",29838 => "0000000000000000",
29839 => "0000000000000000",29840 => "0000000000000000",
29841 => "0000000000000000",29842 => "0000000000000000",
29843 => "0000000000000000",29844 => "0000000000000000",
29845 => "0000000000000000",29846 => "0000000000000000",
29847 => "0000000000000000",29848 => "0000000000000000",
29849 => "0000000000000000",29850 => "0000000000000000",
29851 => "0000000000000000",29852 => "0000000000000000",
29853 => "0000000000000000",29854 => "0000000000000000",
29855 => "0000000000000000",29856 => "0000000000000000",
29857 => "0000000000000000",29858 => "0000000000000000",
29859 => "0000000000000000",29860 => "0000000000000000",
29861 => "0000000000000000",29862 => "0000000000000000",
29863 => "0000000000000000",29864 => "0000000000000000",
29865 => "0000000000000000",29866 => "0000000000000000",
29867 => "0000000000000000",29868 => "0000000000000000",
29869 => "0000000000000000",29870 => "0000000000000000",
29871 => "0000000000000000",29872 => "0000000000000000",
29873 => "0000000000000000",29874 => "0000000000000000",
29875 => "0000000000000000",29876 => "0000000000000000",
29877 => "0000000000000000",29878 => "0000000000000000",
29879 => "0000000000000000",29880 => "0000000000000000",
29881 => "0000000000000000",29882 => "0000000000000000",
29883 => "0000000000000000",29884 => "0000000000000000",
29885 => "0000000000000000",29886 => "0000000000000000",
29887 => "0000000000000000",29888 => "0000000000000000",
29889 => "0000000000000000",29890 => "0000000000000000",
29891 => "0000000000000000",29892 => "0000000000000000",
29893 => "0000000000000000",29894 => "0000000000000000",
29895 => "0000000000000000",29896 => "0000000000000000",
29897 => "0000000000000000",29898 => "0000000000000000",
29899 => "0000000000000000",29900 => "0000000000000000",
29901 => "0000000000000000",29902 => "0000000000000000",
29903 => "0000000000000000",29904 => "0000000000000000",
29905 => "0000000000000000",29906 => "0000000000000000",
29907 => "0000000000000000",29908 => "0000000000000000",
29909 => "0000000000000000",29910 => "0000000000000000",
29911 => "0000000000000000",29912 => "0000000000000000",
29913 => "0000000000000000",29914 => "0000000000000000",
29915 => "0000000000000000",29916 => "0000000000000000",
29917 => "0000000000000000",29918 => "0000000000000000",
29919 => "0000000000000000",29920 => "0000000000000000",
29921 => "0000000000000000",29922 => "0000000000000000",
29923 => "0000000000000000",29924 => "0000000000000000",
29925 => "0000000000000000",29926 => "0000000000000000",
29927 => "0000000000000000",29928 => "0000000000000000",
29929 => "0000000000000000",29930 => "0000000000000000",
29931 => "0000000000000000",29932 => "0000000000000000",
29933 => "0000000000000000",29934 => "0000000000000000",
29935 => "0000000000000000",29936 => "0000000000000000",
29937 => "0000000000000000",29938 => "0000000000000000",
29939 => "0000000000000000",29940 => "0000000000000000",
29941 => "0000000000000000",29942 => "0000000000000000",
29943 => "0000000000000000",29944 => "0000000000000000",
29945 => "0000000000000000",29946 => "0000000000000000",
29947 => "0000000000000000",29948 => "0000000000000000",
29949 => "0000000000000000",29950 => "0000000000000000",
29951 => "0000000000000000",29952 => "0000000000000000",
29953 => "0000000000000000",29954 => "0000000000000000",
29955 => "0000000000000000",29956 => "0000000000000000",
29957 => "0000000000000000",29958 => "0000000000000000",
29959 => "0000000000000000",29960 => "0000000000000000",
29961 => "0000000000000000",29962 => "0000000000000000",
29963 => "0000000000000000",29964 => "0000000000000000",
29965 => "0000000000000000",29966 => "0000000000000000",
29967 => "0000000000000000",29968 => "0000000000000000",
29969 => "0000000000000000",29970 => "0000000000000000",
29971 => "0000000000000000",29972 => "0000000000000000",
29973 => "0000000000000000",29974 => "0000000000000000",
29975 => "0000000000000000",29976 => "0000000000000000",
29977 => "0000000000000000",29978 => "0000000000000000",
29979 => "0000000000000000",29980 => "0000000000000000",
29981 => "0000000000000000",29982 => "0000000000000000",
29983 => "0000000000000000",29984 => "0000000000000000",
29985 => "0000000000000000",29986 => "0000000000000000",
29987 => "0000000000000000",29988 => "0000000000000000",
29989 => "0000000000000000",29990 => "0000000000000000",
29991 => "0000000000000000",29992 => "0000000000000000",
29993 => "0000000000000000",29994 => "0000000000000000",
29995 => "0000000000000000",29996 => "0000000000000000",
29997 => "0000000000000000",29998 => "0000000000000000",
29999 => "0000000000000000",30000 => "0000000000000000",
30001 => "0000000000000000",30002 => "0000000000000000",
30003 => "0000000000000000",30004 => "0000000000000000",
30005 => "0000000000000000",30006 => "0000000000000000",
30007 => "0000000000000000",30008 => "0000000000000000",
30009 => "0000000000000000",30010 => "0000000000000000",
30011 => "0000000000000000",30012 => "0000000000000000",
30013 => "0000000000000000",30014 => "0000000000000000",
30015 => "0000000000000000",30016 => "0000000000000000",
30017 => "0000000000000000",30018 => "0000000000000000",
30019 => "0000000000000000",30020 => "0000000000000000",
30021 => "0000000000000000",30022 => "0000000000000000",
30023 => "0000000000000000",30024 => "0000000000000000",
30025 => "0000000000000000",30026 => "0000000000000000",
30027 => "0000000000000000",30028 => "0000000000000000",
30029 => "0000000000000000",30030 => "0000000000000000",
30031 => "0000000000000000",30032 => "0000000000000000",
30033 => "0000000000000000",30034 => "0000000000000000",
30035 => "0000000000000000",30036 => "0000000000000000",
30037 => "0000000000000000",30038 => "0000000000000000",
30039 => "0000000000000000",30040 => "0000000000000000",
30041 => "0000000000000000",30042 => "0000000000000000",
30043 => "0000000000000000",30044 => "0000000000000000",
30045 => "0000000000000000",30046 => "0000000000000000",
30047 => "0000000000000000",30048 => "0000000000000000",
30049 => "0000000000000000",30050 => "0000000000000000",
30051 => "0000000000000000",30052 => "0000000000000000",
30053 => "0000000000000000",30054 => "0000000000000000",
30055 => "0000000000000000",30056 => "0000000000000000",
30057 => "0000000000000000",30058 => "0000000000000000",
30059 => "0000000000000000",30060 => "0000000000000000",
30061 => "0000000000000000",30062 => "0000000000000000",
30063 => "0000000000000000",30064 => "0000000000000000",
30065 => "0000000000000000",30066 => "0000000000000000",
30067 => "0000000000000000",30068 => "0000000000000000",
30069 => "0000000000000000",30070 => "0000000000000000",
30071 => "0000000000000000",30072 => "0000000000000000",
30073 => "0000000000000000",30074 => "0000000000000000",
30075 => "0000000000000000",30076 => "0000000000000000",
30077 => "0000000000000000",30078 => "0000000000000000",
30079 => "0000000000000000",30080 => "0000000000000000",
30081 => "0000000000000000",30082 => "0000000000000000",
30083 => "0000000000000000",30084 => "0000000000000000",
30085 => "0000000000000000",30086 => "0000000000000000",
30087 => "0000000000000000",30088 => "0000000000000000",
30089 => "0000000000000000",30090 => "0000000000000000",
30091 => "0000000000000000",30092 => "0000000000000000",
30093 => "0000000000000000",30094 => "0000000000000000",
30095 => "0000000000000000",30096 => "0000000000000000",
30097 => "0000000000000000",30098 => "0000000000000000",
30099 => "0000000000000000",30100 => "0000000000000000",
30101 => "0000000000000000",30102 => "0000000000000000",
30103 => "0000000000000000",30104 => "0000000000000000",
30105 => "0000000000000000",30106 => "0000000000000000",
30107 => "0000000000000000",30108 => "0000000000000000",
30109 => "0000000000000000",30110 => "0000000000000000",
30111 => "0000000000000000",30112 => "0000000000000000",
30113 => "0000000000000000",30114 => "0000000000000000",
30115 => "0000000000000000",30116 => "0000000000000000",
30117 => "0000000000000000",30118 => "0000000000000000",
30119 => "0000000000000000",30120 => "0000000000000000",
30121 => "0000000000000000",30122 => "0000000000000000",
30123 => "0000000000000000",30124 => "0000000000000000",
30125 => "0000000000000000",30126 => "0000000000000000",
30127 => "0000000000000000",30128 => "0000000000000000",
30129 => "0000000000000000",30130 => "0000000000000000",
30131 => "0000000000000000",30132 => "0000000000000000",
30133 => "0000000000000000",30134 => "0000000000000000",
30135 => "0000000000000000",30136 => "0000000000000000",
30137 => "0000000000000000",30138 => "0000000000000000",
30139 => "0000000000000000",30140 => "0000000000000000",
30141 => "0000000000000000",30142 => "0000000000000000",
30143 => "0000000000000000",30144 => "0000000000000000",
30145 => "0000000000000000",30146 => "0000000000000000",
30147 => "0000000000000000",30148 => "0000000000000000",
30149 => "0000000000000000",30150 => "0000000000000000",
30151 => "0000000000000000",30152 => "0000000000000000",
30153 => "0000000000000000",30154 => "0000000000000000",
30155 => "0000000000000000",30156 => "0000000000000000",
30157 => "0000000000000000",30158 => "0000000000000000",
30159 => "0000000000000000",30160 => "0000000000000000",
30161 => "0000000000000000",30162 => "0000000000000000",
30163 => "0000000000000000",30164 => "0000000000000000",
30165 => "0000000000000000",30166 => "0000000000000000",
30167 => "0000000000000000",30168 => "0000000000000000",
30169 => "0000000000000000",30170 => "0000000000000000",
30171 => "0000000000000000",30172 => "0000000000000000",
30173 => "0000000000000000",30174 => "0000000000000000",
30175 => "0000000000000000",30176 => "0000000000000000",
30177 => "0000000000000000",30178 => "0000000000000000",
30179 => "0000000000000000",30180 => "0000000000000000",
30181 => "0000000000000000",30182 => "0000000000000000",
30183 => "0000000000000000",30184 => "0000000000000000",
30185 => "0000000000000000",30186 => "0000000000000000",
30187 => "0000000000000000",30188 => "0000000000000000",
30189 => "0000000000000000",30190 => "0000000000000000",
30191 => "0000000000000000",30192 => "0000000000000000",
30193 => "0000000000000000",30194 => "0000000000000000",
30195 => "0000000000000000",30196 => "0000000000000000",
30197 => "0000000000000000",30198 => "0000000000000000",
30199 => "0000000000000000",30200 => "0000000000000000",
30201 => "0000000000000000",30202 => "0000000000000000",
30203 => "0000000000000000",30204 => "0000000000000000",
30205 => "0000000000000000",30206 => "0000000000000000",
30207 => "0000000000000000",30208 => "0000000000000000",
30209 => "0000000000000000",30210 => "0000000000000000",
30211 => "0000000000000000",30212 => "0000000000000000",
30213 => "0000000000000000",30214 => "0000000000000000",
30215 => "0000000000000000",30216 => "0000000000000000",
30217 => "0000000000000000",30218 => "0000000000000000",
30219 => "0000000000000000",30220 => "0000000000000000",
30221 => "0000000000000000",30222 => "0000000000000000",
30223 => "0000000000000000",30224 => "0000000000000000",
30225 => "0000000000000000",30226 => "0000000000000000",
30227 => "0000000000000000",30228 => "0000000000000000",
30229 => "0000000000000000",30230 => "0000000000000000",
30231 => "0000000000000000",30232 => "0000000000000000",
30233 => "0000000000000000",30234 => "0000000000000000",
30235 => "0000000000000000",30236 => "0000000000000000",
30237 => "0000000000000000",30238 => "0000000000000000",
30239 => "0000000000000000",30240 => "0000000000000000",
30241 => "0000000000000000",30242 => "0000000000000000",
30243 => "0000000000000000",30244 => "0000000000000000",
30245 => "0000000000000000",30246 => "0000000000000000",
30247 => "0000000000000000",30248 => "0000000000000000",
30249 => "0000000000000000",30250 => "0000000000000000",
30251 => "0000000000000000",30252 => "0000000000000000",
30253 => "0000000000000000",30254 => "0000000000000000",
30255 => "0000000000000000",30256 => "0000000000000000",
30257 => "0000000000000000",30258 => "0000000000000000",
30259 => "0000000000000000",30260 => "0000000000000000",
30261 => "0000000000000000",30262 => "0000000000000000",
30263 => "0000000000000000",30264 => "0000000000000000",
30265 => "0000000000000000",30266 => "0000000000000000",
30267 => "0000000000000000",30268 => "0000000000000000",
30269 => "0000000000000000",30270 => "0000000000000000",
30271 => "0000000000000000",30272 => "0000000000000000",
30273 => "0000000000000000",30274 => "0000000000000000",
30275 => "0000000000000000",30276 => "0000000000000000",
30277 => "0000000000000000",30278 => "0000000000000000",
30279 => "0000000000000000",30280 => "0000000000000000",
30281 => "0000000000000000",30282 => "0000000000000000",
30283 => "0000000000000000",30284 => "0000000000000000",
30285 => "0000000000000000",30286 => "0000000000000000",
30287 => "0000000000000000",30288 => "0000000000000000",
30289 => "0000000000000000",30290 => "0000000000000000",
30291 => "0000000000000000",30292 => "0000000000000000",
30293 => "0000000000000000",30294 => "0000000000000000",
30295 => "0000000000000000",30296 => "0000000000000000",
30297 => "0000000000000000",30298 => "0000000000000000",
30299 => "0000000000000000",30300 => "0000000000000000",
30301 => "0000000000000000",30302 => "0000000000000000",
30303 => "0000000000000000",30304 => "0000000000000000",
30305 => "0000000000000000",30306 => "0000000000000000",
30307 => "0000000000000000",30308 => "0000000000000000",
30309 => "0000000000000000",30310 => "0000000000000000",
30311 => "0000000000000000",30312 => "0000000000000000",
30313 => "0000000000000000",30314 => "0000000000000000",
30315 => "0000000000000000",30316 => "0000000000000000",
30317 => "0000000000000000",30318 => "0000000000000000",
30319 => "0000000000000000",30320 => "0000000000000000",
30321 => "0000000000000000",30322 => "0000000000000000",
30323 => "0000000000000000",30324 => "0000000000000000",
30325 => "0000000000000000",30326 => "0000000000000000",
30327 => "0000000000000000",30328 => "0000000000000000",
30329 => "0000000000000000",30330 => "0000000000000000",
30331 => "0000000000000000",30332 => "0000000000000000",
30333 => "0000000000000000",30334 => "0000000000000000",
30335 => "0000000000000000",30336 => "0000000000000000",
30337 => "0000000000000000",30338 => "0000000000000000",
30339 => "0000000000000000",30340 => "0000000000000000",
30341 => "0000000000000000",30342 => "0000000000000000",
30343 => "0000000000000000",30344 => "0000000000000000",
30345 => "0000000000000000",30346 => "0000000000000000",
30347 => "0000000000000000",30348 => "0000000000000000",
30349 => "0000000000000000",30350 => "0000000000000000",
30351 => "0000000000000000",30352 => "0000000000000000",
30353 => "0000000000000000",30354 => "0000000000000000",
30355 => "0000000000000000",30356 => "0000000000000000",
30357 => "0000000000000000",30358 => "0000000000000000",
30359 => "0000000000000000",30360 => "0000000000000000",
30361 => "0000000000000000",30362 => "0000000000000000",
30363 => "0000000000000000",30364 => "0000000000000000",
30365 => "0000000000000000",30366 => "0000000000000000",
30367 => "0000000000000000",30368 => "0000000000000000",
30369 => "0000000000000000",30370 => "0000000000000000",
30371 => "0000000000000000",30372 => "0000000000000000",
30373 => "0000000000000000",30374 => "0000000000000000",
30375 => "0000000000000000",30376 => "0000000000000000",
30377 => "0000000000000000",30378 => "0000000000000000",
30379 => "0000000000000000",30380 => "0000000000000000",
30381 => "0000000000000000",30382 => "0000000000000000",
30383 => "0000000000000000",30384 => "0000000000000000",
30385 => "0000000000000000",30386 => "0000000000000000",
30387 => "0000000000000000",30388 => "0000000000000000",
30389 => "0000000000000000",30390 => "0000000000000000",
30391 => "0000000000000000",30392 => "0000000000000000",
30393 => "0000000000000000",30394 => "0000000000000000",
30395 => "0000000000000000",30396 => "0000000000000000",
30397 => "0000000000000000",30398 => "0000000000000000",
30399 => "0000000000000000",30400 => "0000000000000000",
30401 => "0000000000000000",30402 => "0000000000000000",
30403 => "0000000000000000",30404 => "0000000000000000",
30405 => "0000000000000000",30406 => "0000000000000000",
30407 => "0000000000000000",30408 => "0000000000000000",
30409 => "0000000000000000",30410 => "0000000000000000",
30411 => "0000000000000000",30412 => "0000000000000000",
30413 => "0000000000000000",30414 => "0000000000000000",
30415 => "0000000000000000",30416 => "0000000000000000",
30417 => "0000000000000000",30418 => "0000000000000000",
30419 => "0000000000000000",30420 => "0000000000000000",
30421 => "0000000000000000",30422 => "0000000000000000",
30423 => "0000000000000000",30424 => "0000000000000000",
30425 => "0000000000000000",30426 => "0000000000000000",
30427 => "0000000000000000",30428 => "0000000000000000",
30429 => "0000000000000000",30430 => "0000000000000000",
30431 => "0000000000000000",30432 => "0000000000000000",
30433 => "0000000000000000",30434 => "0000000000000000",
30435 => "0000000000000000",30436 => "0000000000000000",
30437 => "0000000000000000",30438 => "0000000000000000",
30439 => "0000000000000000",30440 => "0000000000000000",
30441 => "0000000000000000",30442 => "0000000000000000",
30443 => "0000000000000000",30444 => "0000000000000000",
30445 => "0000000000000000",30446 => "0000000000000000",
30447 => "0000000000000000",30448 => "0000000000000000",
30449 => "0000000000000000",30450 => "0000000000000000",
30451 => "0000000000000000",30452 => "0000000000000000",
30453 => "0000000000000000",30454 => "0000000000000000",
30455 => "0000000000000000",30456 => "0000000000000000",
30457 => "0000000000000000",30458 => "0000000000000000",
30459 => "0000000000000000",30460 => "0000000000000000",
30461 => "0000000000000000",30462 => "0000000000000000",
30463 => "0000000000000000",30464 => "0000000000000000",
30465 => "0000000000000000",30466 => "0000000000000000",
30467 => "0000000000000000",30468 => "0000000000000000",
30469 => "0000000000000000",30470 => "0000000000000000",
30471 => "0000000000000000",30472 => "0000000000000000",
30473 => "0000000000000000",30474 => "0000000000000000",
30475 => "0000000000000000",30476 => "0000000000000000",
30477 => "0000000000000000",30478 => "0000000000000000",
30479 => "0000000000000000",30480 => "0000000000000000",
30481 => "0000000000000000",30482 => "0000000000000000",
30483 => "0000000000000000",30484 => "0000000000000000",
30485 => "0000000000000000",30486 => "0000000000000000",
30487 => "0000000000000000",30488 => "0000000000000000",
30489 => "0000000000000000",30490 => "0000000000000000",
30491 => "0000000000000000",30492 => "0000000000000000",
30493 => "0000000000000000",30494 => "0000000000000000",
30495 => "0000000000000000",30496 => "0000000000000000",
30497 => "0000000000000000",30498 => "0000000000000000",
30499 => "0000000000000000",30500 => "0000000000000000",
30501 => "0000000000000000",30502 => "0000000000000000",
30503 => "0000000000000000",30504 => "0000000000000000",
30505 => "0000000000000000",30506 => "0000000000000000",
30507 => "0000000000000000",30508 => "0000000000000000",
30509 => "0000000000000000",30510 => "0000000000000000",
30511 => "0000000000000000",30512 => "0000000000000000",
30513 => "0000000000000000",30514 => "0000000000000000",
30515 => "0000000000000000",30516 => "0000000000000000",
30517 => "0000000000000000",30518 => "0000000000000000",
30519 => "0000000000000000",30520 => "0000000000000000",
30521 => "0000000000000000",30522 => "0000000000000000",
30523 => "0000000000000000",30524 => "0000000000000000",
30525 => "0000000000000000",30526 => "0000000000000000",
30527 => "0000000000000000",30528 => "0000000000000000",
30529 => "0000000000000000",30530 => "0000000000000000",
30531 => "0000000000000000",30532 => "0000000000000000",
30533 => "0000000000000000",30534 => "0000000000000000",
30535 => "0000000000000000",30536 => "0000000000000000",
30537 => "0000000000000000",30538 => "0000000000000000",
30539 => "0000000000000000",30540 => "0000000000000000",
30541 => "0000000000000000",30542 => "0000000000000000",
30543 => "0000000000000000",30544 => "0000000000000000",
30545 => "0000000000000000",30546 => "0000000000000000",
30547 => "0000000000000000",30548 => "0000000000000000",
30549 => "0000000000000000",30550 => "0000000000000000",
30551 => "0000000000000000",30552 => "0000000000000000",
30553 => "0000000000000000",30554 => "0000000000000000",
30555 => "0000000000000000",30556 => "0000000000000000",
30557 => "0000000000000000",30558 => "0000000000000000",
30559 => "0000000000000000",30560 => "0000000000000000",
30561 => "0000000000000000",30562 => "0000000000000000",
30563 => "0000000000000000",30564 => "0000000000000000",
30565 => "0000000000000000",30566 => "0000000000000000",
30567 => "0000000000000000",30568 => "0000000000000000",
30569 => "0000000000000000",30570 => "0000000000000000",
30571 => "0000000000000000",30572 => "0000000000000000",
30573 => "0000000000000000",30574 => "0000000000000000",
30575 => "0000000000000000",30576 => "0000000000000000",
30577 => "0000000000000000",30578 => "0000000000000000",
30579 => "0000000000000000",30580 => "0000000000000000",
30581 => "0000000000000000",30582 => "0000000000000000",
30583 => "0000000000000000",30584 => "0000000000000000",
30585 => "0000000000000000",30586 => "0000000000000000",
30587 => "0000000000000000",30588 => "0000000000000000",
30589 => "0000000000000000",30590 => "0000000000000000",
30591 => "0000000000000000",30592 => "0000000000000000",
30593 => "0000000000000000",30594 => "0000000000000000",
30595 => "0000000000000000",30596 => "0000000000000000",
30597 => "0000000000000000",30598 => "0000000000000000",
30599 => "0000000000000000",30600 => "0000000000000000",
30601 => "0000000000000000",30602 => "0000000000000000",
30603 => "0000000000000000",30604 => "0000000000000000",
30605 => "0000000000000000",30606 => "0000000000000000",
30607 => "0000000000000000",30608 => "0000000000000000",
30609 => "0000000000000000",30610 => "0000000000000000",
30611 => "0000000000000000",30612 => "0000000000000000",
30613 => "0000000000000000",30614 => "0000000000000000",
30615 => "0000000000000000",30616 => "0000000000000000",
30617 => "0000000000000000",30618 => "0000000000000000",
30619 => "0000000000000000",30620 => "0000000000000000",
30621 => "0000000000000000",30622 => "0000000000000000",
30623 => "0000000000000000",30624 => "0000000000000000",
30625 => "0000000000000000",30626 => "0000000000000000",
30627 => "0000000000000000",30628 => "0000000000000000",
30629 => "0000000000000000",30630 => "0000000000000000",
30631 => "0000000000000000",30632 => "0000000000000000",
30633 => "0000000000000000",30634 => "0000000000000000",
30635 => "0000000000000000",30636 => "0000000000000000",
30637 => "0000000000000000",30638 => "0000000000000000",
30639 => "0000000000000000",30640 => "0000000000000000",
30641 => "0000000000000000",30642 => "0000000000000000",
30643 => "0000000000000000",30644 => "0000000000000000",
30645 => "0000000000000000",30646 => "0000000000000000",
30647 => "0000000000000000",30648 => "0000000000000000",
30649 => "0000000000000000",30650 => "0000000000000000",
30651 => "0000000000000000",30652 => "0000000000000000",
30653 => "0000000000000000",30654 => "0000000000000000",
30655 => "0000000000000000",30656 => "0000000000000000",
30657 => "0000000000000000",30658 => "0000000000000000",
30659 => "0000000000000000",30660 => "0000000000000000",
30661 => "0000000000000000",30662 => "0000000000000000",
30663 => "0000000000000000",30664 => "0000000000000000",
30665 => "0000000000000000",30666 => "0000000000000000",
30667 => "0000000000000000",30668 => "0000000000000000",
30669 => "0000000000000000",30670 => "0000000000000000",
30671 => "0000000000000000",30672 => "0000000000000000",
30673 => "0000000000000000",30674 => "0000000000000000",
30675 => "0000000000000000",30676 => "0000000000000000",
30677 => "0000000000000000",30678 => "0000000000000000",
30679 => "0000000000000000",30680 => "0000000000000000",
30681 => "0000000000000000",30682 => "0000000000000000",
30683 => "0000000000000000",30684 => "0000000000000000",
30685 => "0000000000000000",30686 => "0000000000000000",
30687 => "0000000000000000",30688 => "0000000000000000",
30689 => "0000000000000000",30690 => "0000000000000000",
30691 => "0000000000000000",30692 => "0000000000000000",
30693 => "0000000000000000",30694 => "0000000000000000",
30695 => "0000000000000000",30696 => "0000000000000000",
30697 => "0000000000000000",30698 => "0000000000000000",
30699 => "0000000000000000",30700 => "0000000000000000",
30701 => "0000000000000000",30702 => "0000000000000000",
30703 => "0000000000000000",30704 => "0000000000000000",
30705 => "0000000000000000",30706 => "0000000000000000",
30707 => "0000000000000000",30708 => "0000000000000000",
30709 => "0000000000000000",30710 => "0000000000000000",
30711 => "0000000000000000",30712 => "0000000000000000",
30713 => "0000000000000000",30714 => "0000000000000000",
30715 => "0000000000000000",30716 => "0000000000000000",
30717 => "0000000000000000",30718 => "0000000000000000",
30719 => "0000000000000000",30720 => "0000000000000000",
30721 => "0000000000000000",30722 => "0000000000000000",
30723 => "0000000000000000",30724 => "0000000000000000",
30725 => "0000000000000000",30726 => "0000000000000000",
30727 => "0000000000000000",30728 => "0000000000000000",
30729 => "0000000000000000",30730 => "0000000000000000",
30731 => "0000000000000000",30732 => "0000000000000000",
30733 => "0000000000000000",30734 => "0000000000000000",
30735 => "0000000000000000",30736 => "0000000000000000",
30737 => "0000000000000000",30738 => "0000000000000000",
30739 => "0000000000000000",30740 => "0000000000000000",
30741 => "0000000000000000",30742 => "0000000000000000",
30743 => "0000000000000000",30744 => "0000000000000000",
30745 => "0000000000000000",30746 => "0000000000000000",
30747 => "0000000000000000",30748 => "0000000000000000",
30749 => "0000000000000000",30750 => "0000000000000000",
30751 => "0000000000000000",30752 => "0000000000000000",
30753 => "0000000000000000",30754 => "0000000000000000",
30755 => "0000000000000000",30756 => "0000000000000000",
30757 => "0000000000000000",30758 => "0000000000000000",
30759 => "0000000000000000",30760 => "0000000000000000",
30761 => "0000000000000000",30762 => "0000000000000000",
30763 => "0000000000000000",30764 => "0000000000000000",
30765 => "0000000000000000",30766 => "0000000000000000",
30767 => "0000000000000000",30768 => "0000000000000000",
30769 => "0000000000000000",30770 => "0000000000000000",
30771 => "0000000000000000",30772 => "0000000000000000",
30773 => "0000000000000000",30774 => "0000000000000000",
30775 => "0000000000000000",30776 => "0000000000000000",
30777 => "0000000000000000",30778 => "0000000000000000",
30779 => "0000000000000000",30780 => "0000000000000000",
30781 => "0000000000000000",30782 => "0000000000000000",
30783 => "0000000000000000",30784 => "0000000000000000",
30785 => "0000000000000000",30786 => "0000000000000000",
30787 => "0000000000000000",30788 => "0000000000000000",
30789 => "0000000000000000",30790 => "0000000000000000",
30791 => "0000000000000000",30792 => "0000000000000000",
30793 => "0000000000000000",30794 => "0000000000000000",
30795 => "0000000000000000",30796 => "0000000000000000",
30797 => "0000000000000000",30798 => "0000000000000000",
30799 => "0000000000000000",30800 => "0000000000000000",
30801 => "0000000000000000",30802 => "0000000000000000",
30803 => "0000000000000000",30804 => "0000000000000000",
30805 => "0000000000000000",30806 => "0000000000000000",
30807 => "0000000000000000",30808 => "0000000000000000",
30809 => "0000000000000000",30810 => "0000000000000000",
30811 => "0000000000000000",30812 => "0000000000000000",
30813 => "0000000000000000",30814 => "0000000000000000",
30815 => "0000000000000000",30816 => "0000000000000000",
30817 => "0000000000000000",30818 => "0000000000000000",
30819 => "0000000000000000",30820 => "0000000000000000",
30821 => "0000000000000000",30822 => "0000000000000000",
30823 => "0000000000000000",30824 => "0000000000000000",
30825 => "0000000000000000",30826 => "0000000000000000",
30827 => "0000000000000000",30828 => "0000000000000000",
30829 => "0000000000000000",30830 => "0000000000000000",
30831 => "0000000000000000",30832 => "0000000000000000",
30833 => "0000000000000000",30834 => "0000000000000000",
30835 => "0000000000000000",30836 => "0000000000000000",
30837 => "0000000000000000",30838 => "0000000000000000",
30839 => "0000000000000000",30840 => "0000000000000000",
30841 => "0000000000000000",30842 => "0000000000000000",
30843 => "0000000000000000",30844 => "0000000000000000",
30845 => "0000000000000000",30846 => "0000000000000000",
30847 => "0000000000000000",30848 => "0000000000000000",
30849 => "0000000000000000",30850 => "0000000000000000",
30851 => "0000000000000000",30852 => "0000000000000000",
30853 => "0000000000000000",30854 => "0000000000000000",
30855 => "0000000000000000",30856 => "0000000000000000",
30857 => "0000000000000000",30858 => "0000000000000000",
30859 => "0000000000000000",30860 => "0000000000000000",
30861 => "0000000000000000",30862 => "0000000000000000",
30863 => "0000000000000000",30864 => "0000000000000000",
30865 => "0000000000000000",30866 => "0000000000000000",
30867 => "0000000000000000",30868 => "0000000000000000",
30869 => "0000000000000000",30870 => "0000000000000000",
30871 => "0000000000000000",30872 => "0000000000000000",
30873 => "0000000000000000",30874 => "0000000000000000",
30875 => "0000000000000000",30876 => "0000000000000000",
30877 => "0000000000000000",30878 => "0000000000000000",
30879 => "0000000000000000",30880 => "0000000000000000",
30881 => "0000000000000000",30882 => "0000000000000000",
30883 => "0000000000000000",30884 => "0000000000000000",
30885 => "0000000000000000",30886 => "0000000000000000",
30887 => "0000000000000000",30888 => "0000000000000000",
30889 => "0000000000000000",30890 => "0000000000000000",
30891 => "0000000000000000",30892 => "0000000000000000",
30893 => "0000000000000000",30894 => "0000000000000000",
30895 => "0000000000000000",30896 => "0000000000000000",
30897 => "0000000000000000",30898 => "0000000000000000",
30899 => "0000000000000000",30900 => "0000000000000000",
30901 => "0000000000000000",30902 => "0000000000000000",
30903 => "0000000000000000",30904 => "0000000000000000",
30905 => "0000000000000000",30906 => "0000000000000000",
30907 => "0000000000000000",30908 => "0000000000000000",
30909 => "0000000000000000",30910 => "0000000000000000",
30911 => "0000000000000000",30912 => "0000000000000000",
30913 => "0000000000000000",30914 => "0000000000000000",
30915 => "0000000000000000",30916 => "0000000000000000",
30917 => "0000000000000000",30918 => "0000000000000000",
30919 => "0000000000000000",30920 => "0000000000000000",
30921 => "0000000000000000",30922 => "0000000000000000",
30923 => "0000000000000000",30924 => "0000000000000000",
30925 => "0000000000000000",30926 => "0000000000000000",
30927 => "0000000000000000",30928 => "0000000000000000",
30929 => "0000000000000000",30930 => "0000000000000000",
30931 => "0000000000000000",30932 => "0000000000000000",
30933 => "0000000000000000",30934 => "0000000000000000",
30935 => "0000000000000000",30936 => "0000000000000000",
30937 => "0000000000000000",30938 => "0000000000000000",
30939 => "0000000000000000",30940 => "0000000000000000",
30941 => "0000000000000000",30942 => "0000000000000000",
30943 => "0000000000000000",30944 => "0000000000000000",
30945 => "0000000000000000",30946 => "0000000000000000",
30947 => "0000000000000000",30948 => "0000000000000000",
30949 => "0000000000000000",30950 => "0000000000000000",
30951 => "0000000000000000",30952 => "0000000000000000",
30953 => "0000000000000000",30954 => "0000000000000000",
30955 => "0000000000000000",30956 => "0000000000000000",
30957 => "0000000000000000",30958 => "0000000000000000",
30959 => "0000000000000000",30960 => "0000000000000000",
30961 => "0000000000000000",30962 => "0000000000000000",
30963 => "0000000000000000",30964 => "0000000000000000",
30965 => "0000000000000000",30966 => "0000000000000000",
30967 => "0000000000000000",30968 => "0000000000000000",
30969 => "0000000000000000",30970 => "0000000000000000",
30971 => "0000000000000000",30972 => "0000000000000000",
30973 => "0000000000000000",30974 => "0000000000000000",
30975 => "0000000000000000",30976 => "0000000000000000",
30977 => "0000000000000000",30978 => "0000000000000000",
30979 => "0000000000000000",30980 => "0000000000000000",
30981 => "0000000000000000",30982 => "0000000000000000",
30983 => "0000000000000000",30984 => "0000000000000000",
30985 => "0000000000000000",30986 => "0000000000000000",
30987 => "0000000000000000",30988 => "0000000000000000",
30989 => "0000000000000000",30990 => "0000000000000000",
30991 => "0000000000000000",30992 => "0000000000000000",
30993 => "0000000000000000",30994 => "0000000000000000",
30995 => "0000000000000000",30996 => "0000000000000000",
30997 => "0000000000000000",30998 => "0000000000000000",
30999 => "0000000000000000",31000 => "0000000000000000",
31001 => "0000000000000000",31002 => "0000000000000000",
31003 => "0000000000000000",31004 => "0000000000000000",
31005 => "0000000000000000",31006 => "0000000000000000",
31007 => "0000000000000000",31008 => "0000000000000000",
31009 => "0000000000000000",31010 => "0000000000000000",
31011 => "0000000000000000",31012 => "0000000000000000",
31013 => "0000000000000000",31014 => "0000000000000000",
31015 => "0000000000000000",31016 => "0000000000000000",
31017 => "0000000000000000",31018 => "0000000000000000",
31019 => "0000000000000000",31020 => "0000000000000000",
31021 => "0000000000000000",31022 => "0000000000000000",
31023 => "0000000000000000",31024 => "0000000000000000",
31025 => "0000000000000000",31026 => "0000000000000000",
31027 => "0000000000000000",31028 => "0000000000000000",
31029 => "0000000000000000",31030 => "0000000000000000",
31031 => "0000000000000000",31032 => "0000000000000000",
31033 => "0000000000000000",31034 => "0000000000000000",
31035 => "0000000000000000",31036 => "0000000000000000",
31037 => "0000000000000000",31038 => "0000000000000000",
31039 => "0000000000000000",31040 => "0000000000000000",
31041 => "0000000000000000",31042 => "0000000000000000",
31043 => "0000000000000000",31044 => "0000000000000000",
31045 => "0000000000000000",31046 => "0000000000000000",
31047 => "0000000000000000",31048 => "0000000000000000",
31049 => "0000000000000000",31050 => "0000000000000000",
31051 => "0000000000000000",31052 => "0000000000000000",
31053 => "0000000000000000",31054 => "0000000000000000",
31055 => "0000000000000000",31056 => "0000000000000000",
31057 => "0000000000000000",31058 => "0000000000000000",
31059 => "0000000000000000",31060 => "0000000000000000",
31061 => "0000000000000000",31062 => "0000000000000000",
31063 => "0000000000000000",31064 => "0000000000000000",
31065 => "0000000000000000",31066 => "0000000000000000",
31067 => "0000000000000000",31068 => "0000000000000000",
31069 => "0000000000000000",31070 => "0000000000000000",
31071 => "0000000000000000",31072 => "0000000000000000",
31073 => "0000000000000000",31074 => "0000000000000000",
31075 => "0000000000000000",31076 => "0000000000000000",
31077 => "0000000000000000",31078 => "0000000000000000",
31079 => "0000000000000000",31080 => "0000000000000000",
31081 => "0000000000000000",31082 => "0000000000000000",
31083 => "0000000000000000",31084 => "0000000000000000",
31085 => "0000000000000000",31086 => "0000000000000000",
31087 => "0000000000000000",31088 => "0000000000000000",
31089 => "0000000000000000",31090 => "0000000000000000",
31091 => "0000000000000000",31092 => "0000000000000000",
31093 => "0000000000000000",31094 => "0000000000000000",
31095 => "0000000000000000",31096 => "0000000000000000",
31097 => "0000000000000000",31098 => "0000000000000000",
31099 => "0000000000000000",31100 => "0000000000000000",
31101 => "0000000000000000",31102 => "0000000000000000",
31103 => "0000000000000000",31104 => "0000000000000000",
31105 => "0000000000000000",31106 => "0000000000000000",
31107 => "0000000000000000",31108 => "0000000000000000",
31109 => "0000000000000000",31110 => "0000000000000000",
31111 => "0000000000000000",31112 => "0000000000000000",
31113 => "0000000000000000",31114 => "0000000000000000",
31115 => "0000000000000000",31116 => "0000000000000000",
31117 => "0000000000000000",31118 => "0000000000000000",
31119 => "0000000000000000",31120 => "0000000000000000",
31121 => "0000000000000000",31122 => "0000000000000000",
31123 => "0000000000000000",31124 => "0000000000000000",
31125 => "0000000000000000",31126 => "0000000000000000",
31127 => "0000000000000000",31128 => "0000000000000000",
31129 => "0000000000000000",31130 => "0000000000000000",
31131 => "0000000000000000",31132 => "0000000000000000",
31133 => "0000000000000000",31134 => "0000000000000000",
31135 => "0000000000000000",31136 => "0000000000000000",
31137 => "0000000000000000",31138 => "0000000000000000",
31139 => "0000000000000000",31140 => "0000000000000000",
31141 => "0000000000000000",31142 => "0000000000000000",
31143 => "0000000000000000",31144 => "0000000000000000",
31145 => "0000000000000000",31146 => "0000000000000000",
31147 => "0000000000000000",31148 => "0000000000000000",
31149 => "0000000000000000",31150 => "0000000000000000",
31151 => "0000000000000000",31152 => "0000000000000000",
31153 => "0000000000000000",31154 => "0000000000000000",
31155 => "0000000000000000",31156 => "0000000000000000",
31157 => "0000000000000000",31158 => "0000000000000000",
31159 => "0000000000000000",31160 => "0000000000000000",
31161 => "0000000000000000",31162 => "0000000000000000",
31163 => "0000000000000000",31164 => "0000000000000000",
31165 => "0000000000000000",31166 => "0000000000000000",
31167 => "0000000000000000",31168 => "0000000000000000",
31169 => "0000000000000000",31170 => "0000000000000000",
31171 => "0000000000000000",31172 => "0000000000000000",
31173 => "0000000000000000",31174 => "0000000000000000",
31175 => "0000000000000000",31176 => "0000000000000000",
31177 => "0000000000000000",31178 => "0000000000000000",
31179 => "0000000000000000",31180 => "0000000000000000",
31181 => "0000000000000000",31182 => "0000000000000000",
31183 => "0000000000000000",31184 => "0000000000000000",
31185 => "0000000000000000",31186 => "0000000000000000",
31187 => "0000000000000000",31188 => "0000000000000000",
31189 => "0000000000000000",31190 => "0000000000000000",
31191 => "0000000000000000",31192 => "0000000000000000",
31193 => "0000000000000000",31194 => "0000000000000000",
31195 => "0000000000000000",31196 => "0000000000000000",
31197 => "0000000000000000",31198 => "0000000000000000",
31199 => "0000000000000000",31200 => "0000000000000000",
31201 => "0000000000000000",31202 => "0000000000000000",
31203 => "0000000000000000",31204 => "0000000000000000",
31205 => "0000000000000000",31206 => "0000000000000000",
31207 => "0000000000000000",31208 => "0000000000000000",
31209 => "0000000000000000",31210 => "0000000000000000",
31211 => "0000000000000000",31212 => "0000000000000000",
31213 => "0000000000000000",31214 => "0000000000000000",
31215 => "0000000000000000",31216 => "0000000000000000",
31217 => "0000000000000000",31218 => "0000000000000000",
31219 => "0000000000000000",31220 => "0000000000000000",
31221 => "0000000000000000",31222 => "0000000000000000",
31223 => "0000000000000000",31224 => "0000000000000000",
31225 => "0000000000000000",31226 => "0000000000000000",
31227 => "0000000000000000",31228 => "0000000000000000",
31229 => "0000000000000000",31230 => "0000000000000000",
31231 => "0000000000000000",31232 => "0000000000000000",
31233 => "0000000000000000",31234 => "0000000000000000",
31235 => "0000000000000000",31236 => "0000000000000000",
31237 => "0000000000000000",31238 => "0000000000000000",
31239 => "0000000000000000",31240 => "0000000000000000",
31241 => "0000000000000000",31242 => "0000000000000000",
31243 => "0000000000000000",31244 => "0000000000000000",
31245 => "0000000000000000",31246 => "0000000000000000",
31247 => "0000000000000000",31248 => "0000000000000000",
31249 => "0000000000000000",31250 => "0000000000000000",
31251 => "0000000000000000",31252 => "0000000000000000",
31253 => "0000000000000000",31254 => "0000000000000000",
31255 => "0000000000000000",31256 => "0000000000000000",
31257 => "0000000000000000",31258 => "0000000000000000",
31259 => "0000000000000000",31260 => "0000000000000000",
31261 => "0000000000000000",31262 => "0000000000000000",
31263 => "0000000000000000",31264 => "0000000000000000",
31265 => "0000000000000000",31266 => "0000000000000000",
31267 => "0000000000000000",31268 => "0000000000000000",
31269 => "0000000000000000",31270 => "0000000000000000",
31271 => "0000000000000000",31272 => "0000000000000000",
31273 => "0000000000000000",31274 => "0000000000000000",
31275 => "0000000000000000",31276 => "0000000000000000",
31277 => "0000000000000000",31278 => "0000000000000000",
31279 => "0000000000000000",31280 => "0000000000000000",
31281 => "0000000000000000",31282 => "0000000000000000",
31283 => "0000000000000000",31284 => "0000000000000000",
31285 => "0000000000000000",31286 => "0000000000000000",
31287 => "0000000000000000",31288 => "0000000000000000",
31289 => "0000000000000000",31290 => "0000000000000000",
31291 => "0000000000000000",31292 => "0000000000000000",
31293 => "0000000000000000",31294 => "0000000000000000",
31295 => "0000000000000000",31296 => "0000000000000000",
31297 => "0000000000000000",31298 => "0000000000000000",
31299 => "0000000000000000",31300 => "0000000000000000",
31301 => "0000000000000000",31302 => "0000000000000000",
31303 => "0000000000000000",31304 => "0000000000000000",
31305 => "0000000000000000",31306 => "0000000000000000",
31307 => "0000000000000000",31308 => "0000000000000000",
31309 => "0000000000000000",31310 => "0000000000000000",
31311 => "0000000000000000",31312 => "0000000000000000",
31313 => "0000000000000000",31314 => "0000000000000000",
31315 => "0000000000000000",31316 => "0000000000000000",
31317 => "0000000000000000",31318 => "0000000000000000",
31319 => "0000000000000000",31320 => "0000000000000000",
31321 => "0000000000000000",31322 => "0000000000000000",
31323 => "0000000000000000",31324 => "0000000000000000",
31325 => "0000000000000000",31326 => "0000000000000000",
31327 => "0000000000000000",31328 => "0000000000000000",
31329 => "0000000000000000",31330 => "0000000000000000",
31331 => "0000000000000000",31332 => "0000000000000000",
31333 => "0000000000000000",31334 => "0000000000000000",
31335 => "0000000000000000",31336 => "0000000000000000",
31337 => "0000000000000000",31338 => "0000000000000000",
31339 => "0000000000000000",31340 => "0000000000000000",
31341 => "0000000000000000",31342 => "0000000000000000",
31343 => "0000000000000000",31344 => "0000000000000000",
31345 => "0000000000000000",31346 => "0000000000000000",
31347 => "0000000000000000",31348 => "0000000000000000",
31349 => "0000000000000000",31350 => "0000000000000000",
31351 => "0000000000000000",31352 => "0000000000000000",
31353 => "0000000000000000",31354 => "0000000000000000",
31355 => "0000000000000000",31356 => "0000000000000000",
31357 => "0000000000000000",31358 => "0000000000000000",
31359 => "0000000000000000",31360 => "0000000000000000",
31361 => "0000000000000000",31362 => "0000000000000000",
31363 => "0000000000000000",31364 => "0000000000000000",
31365 => "0000000000000000",31366 => "0000000000000000",
31367 => "0000000000000000",31368 => "0000000000000000",
31369 => "0000000000000000",31370 => "0000000000000000",
31371 => "0000000000000000",31372 => "0000000000000000",
31373 => "0000000000000000",31374 => "0000000000000000",
31375 => "0000000000000000",31376 => "0000000000000000",
31377 => "0000000000000000",31378 => "0000000000000000",
31379 => "0000000000000000",31380 => "0000000000000000",
31381 => "0000000000000000",31382 => "0000000000000000",
31383 => "0000000000000000",31384 => "0000000000000000",
31385 => "0000000000000000",31386 => "0000000000000000",
31387 => "0000000000000000",31388 => "0000000000000000",
31389 => "0000000000000000",31390 => "0000000000000000",
31391 => "0000000000000000",31392 => "0000000000000000",
31393 => "0000000000000000",31394 => "0000000000000000",
31395 => "0000000000000000",31396 => "0000000000000000",
31397 => "0000000000000000",31398 => "0000000000000000",
31399 => "0000000000000000",31400 => "0000000000000000",
31401 => "0000000000000000",31402 => "0000000000000000",
31403 => "0000000000000000",31404 => "0000000000000000",
31405 => "0000000000000000",31406 => "0000000000000000",
31407 => "0000000000000000",31408 => "0000000000000000",
31409 => "0000000000000000",31410 => "0000000000000000",
31411 => "0000000000000000",31412 => "0000000000000000",
31413 => "0000000000000000",31414 => "0000000000000000",
31415 => "0000000000000000",31416 => "0000000000000000",
31417 => "0000000000000000",31418 => "0000000000000000",
31419 => "0000000000000000",31420 => "0000000000000000",
31421 => "0000000000000000",31422 => "0000000000000000",
31423 => "0000000000000000",31424 => "0000000000000000",
31425 => "0000000000000000",31426 => "0000000000000000",
31427 => "0000000000000000",31428 => "0000000000000000",
31429 => "0000000000000000",31430 => "0000000000000000",
31431 => "0000000000000000",31432 => "0000000000000000",
31433 => "0000000000000000",31434 => "0000000000000000",
31435 => "0000000000000000",31436 => "0000000000000000",
31437 => "0000000000000000",31438 => "0000000000000000",
31439 => "0000000000000000",31440 => "0000000000000000",
31441 => "0000000000000000",31442 => "0000000000000000",
31443 => "0000000000000000",31444 => "0000000000000000",
31445 => "0000000000000000",31446 => "0000000000000000",
31447 => "0000000000000000",31448 => "0000000000000000",
31449 => "0000000000000000",31450 => "0000000000000000",
31451 => "0000000000000000",31452 => "0000000000000000",
31453 => "0000000000000000",31454 => "0000000000000000",
31455 => "0000000000000000",31456 => "0000000000000000",
31457 => "0000000000000000",31458 => "0000000000000000",
31459 => "0000000000000000",31460 => "0000000000000000",
31461 => "0000000000000000",31462 => "0000000000000000",
31463 => "0000000000000000",31464 => "0000000000000000",
31465 => "0000000000000000",31466 => "0000000000000000",
31467 => "0000000000000000",31468 => "0000000000000000",
31469 => "0000000000000000",31470 => "0000000000000000",
31471 => "0000000000000000",31472 => "0000000000000000",
31473 => "0000000000000000",31474 => "0000000000000000",
31475 => "0000000000000000",31476 => "0000000000000000",
31477 => "0000000000000000",31478 => "0000000000000000",
31479 => "0000000000000000",31480 => "0000000000000000",
31481 => "0000000000000000",31482 => "0000000000000000",
31483 => "0000000000000000",31484 => "0000000000000000",
31485 => "0000000000000000",31486 => "0000000000000000",
31487 => "0000000000000000",31488 => "0000000000000000",
31489 => "0000000000000000",31490 => "0000000000000000",
31491 => "0000000000000000",31492 => "0000000000000000",
31493 => "0000000000000000",31494 => "0000000000000000",
31495 => "0000000000000000",31496 => "0000000000000000",
31497 => "0000000000000000",31498 => "0000000000000000",
31499 => "0000000000000000",31500 => "0000000000000000",
31501 => "0000000000000000",31502 => "0000000000000000",
31503 => "0000000000000000",31504 => "0000000000000000",
31505 => "0000000000000000",31506 => "0000000000000000",
31507 => "0000000000000000",31508 => "0000000000000000",
31509 => "0000000000000000",31510 => "0000000000000000",
31511 => "0000000000000000",31512 => "0000000000000000",
31513 => "0000000000000000",31514 => "0000000000000000",
31515 => "0000000000000000",31516 => "0000000000000000",
31517 => "0000000000000000",31518 => "0000000000000000",
31519 => "0000000000000000",31520 => "0000000000000000",
31521 => "0000000000000000",31522 => "0000000000000000",
31523 => "0000000000000000",31524 => "0000000000000000",
31525 => "0000000000000000",31526 => "0000000000000000",
31527 => "0000000000000000",31528 => "0000000000000000",
31529 => "0000000000000000",31530 => "0000000000000000",
31531 => "0000000000000000",31532 => "0000000000000000",
31533 => "0000000000000000",31534 => "0000000000000000",
31535 => "0000000000000000",31536 => "0000000000000000",
31537 => "0000000000000000",31538 => "0000000000000000",
31539 => "0000000000000000",31540 => "0000000000000000",
31541 => "0000000000000000",31542 => "0000000000000000",
31543 => "0000000000000000",31544 => "0000000000000000",
31545 => "0000000000000000",31546 => "0000000000000000",
31547 => "0000000000000000",31548 => "0000000000000000",
31549 => "0000000000000000",31550 => "0000000000000000",
31551 => "0000000000000000",31552 => "0000000000000000",
31553 => "0000000000000000",31554 => "0000000000000000",
31555 => "0000000000000000",31556 => "0000000000000000",
31557 => "0000000000000000",31558 => "0000000000000000",
31559 => "0000000000000000",31560 => "0000000000000000",
31561 => "0000000000000000",31562 => "0000000000000000",
31563 => "0000000000000000",31564 => "0000000000000000",
31565 => "0000000000000000",31566 => "0000000000000000",
31567 => "0000000000000000",31568 => "0000000000000000",
31569 => "0000000000000000",31570 => "0000000000000000",
31571 => "0000000000000000",31572 => "0000000000000000",
31573 => "0000000000000000",31574 => "0000000000000000",
31575 => "0000000000000000",31576 => "0000000000000000",
31577 => "0000000000000000",31578 => "0000000000000000",
31579 => "0000000000000000",31580 => "0000000000000000",
31581 => "0000000000000000",31582 => "0000000000000000",
31583 => "0000000000000000",31584 => "0000000000000000",
31585 => "0000000000000000",31586 => "0000000000000000",
31587 => "0000000000000000",31588 => "0000000000000000",
31589 => "0000000000000000",31590 => "0000000000000000",
31591 => "0000000000000000",31592 => "0000000000000000",
31593 => "0000000000000000",31594 => "0000000000000000",
31595 => "0000000000000000",31596 => "0000000000000000",
31597 => "0000000000000000",31598 => "0000000000000000",
31599 => "0000000000000000",31600 => "0000000000000000",
31601 => "0000000000000000",31602 => "0000000000000000",
31603 => "0000000000000000",31604 => "0000000000000000",
31605 => "0000000000000000",31606 => "0000000000000000",
31607 => "0000000000000000",31608 => "0000000000000000",
31609 => "0000000000000000",31610 => "0000000000000000",
31611 => "0000000000000000",31612 => "0000000000000000",
31613 => "0000000000000000",31614 => "0000000000000000",
31615 => "0000000000000000",31616 => "0000000000000000",
31617 => "0000000000000000",31618 => "0000000000000000",
31619 => "0000000000000000",31620 => "0000000000000000",
31621 => "0000000000000000",31622 => "0000000000000000",
31623 => "0000000000000000",31624 => "0000000000000000",
31625 => "0000000000000000",31626 => "0000000000000000",
31627 => "0000000000000000",31628 => "0000000000000000",
31629 => "0000000000000000",31630 => "0000000000000000",
31631 => "0000000000000000",31632 => "0000000000000000",
31633 => "0000000000000000",31634 => "0000000000000000",
31635 => "0000000000000000",31636 => "0000000000000000",
31637 => "0000000000000000",31638 => "0000000000000000",
31639 => "0000000000000000",31640 => "0000000000000000",
31641 => "0000000000000000",31642 => "0000000000000000",
31643 => "0000000000000000",31644 => "0000000000000000",
31645 => "0000000000000000",31646 => "0000000000000000",
31647 => "0000000000000000",31648 => "0000000000000000",
31649 => "0000000000000000",31650 => "0000000000000000",
31651 => "0000000000000000",31652 => "0000000000000000",
31653 => "0000000000000000",31654 => "0000000000000000",
31655 => "0000000000000000",31656 => "0000000000000000",
31657 => "0000000000000000",31658 => "0000000000000000",
31659 => "0000000000000000",31660 => "0000000000000000",
31661 => "0000000000000000",31662 => "0000000000000000",
31663 => "0000000000000000",31664 => "0000000000000000",
31665 => "0000000000000000",31666 => "0000000000000000",
31667 => "0000000000000000",31668 => "0000000000000000",
31669 => "0000000000000000",31670 => "0000000000000000",
31671 => "0000000000000000",31672 => "0000000000000000",
31673 => "0000000000000000",31674 => "0000000000000000",
31675 => "0000000000000000",31676 => "0000000000000000",
31677 => "0000000000000000",31678 => "0000000000000000",
31679 => "0000000000000000",31680 => "0000000000000000",
31681 => "0000000000000000",31682 => "0000000000000000",
31683 => "0000000000000000",31684 => "0000000000000000",
31685 => "0000000000000000",31686 => "0000000000000000",
31687 => "0000000000000000",31688 => "0000000000000000",
31689 => "0000000000000000",31690 => "0000000000000000",
31691 => "0000000000000000",31692 => "0000000000000000",
31693 => "0000000000000000",31694 => "0000000000000000",
31695 => "0000000000000000",31696 => "0000000000000000",
31697 => "0000000000000000",31698 => "0000000000000000",
31699 => "0000000000000000",31700 => "0000000000000000",
31701 => "0000000000000000",31702 => "0000000000000000",
31703 => "0000000000000000",31704 => "0000000000000000",
31705 => "0000000000000000",31706 => "0000000000000000",
31707 => "0000000000000000",31708 => "0000000000000000",
31709 => "0000000000000000",31710 => "0000000000000000",
31711 => "0000000000000000",31712 => "0000000000000000",
31713 => "0000000000000000",31714 => "0000000000000000",
31715 => "0000000000000000",31716 => "0000000000000000",
31717 => "0000000000000000",31718 => "0000000000000000",
31719 => "0000000000000000",31720 => "0000000000000000",
31721 => "0000000000000000",31722 => "0000000000000000",
31723 => "0000000000000000",31724 => "0000000000000000",
31725 => "0000000000000000",31726 => "0000000000000000",
31727 => "0000000000000000",31728 => "0000000000000000",
31729 => "0000000000000000",31730 => "0000000000000000",
31731 => "0000000000000000",31732 => "0000000000000000",
31733 => "0000000000000000",31734 => "0000000000000000",
31735 => "0000000000000000",31736 => "0000000000000000",
31737 => "0000000000000000",31738 => "0000000000000000",
31739 => "0000000000000000",31740 => "0000000000000000",
31741 => "0000000000000000",31742 => "0000000000000000",
31743 => "0000000000000000",31744 => "0000000000000000",
31745 => "0000000000000000",31746 => "0000000000000000",
31747 => "0000000000000000",31748 => "0000000000000000",
31749 => "0000000000000000",31750 => "0000000000000000",
31751 => "0000000000000000",31752 => "0000000000000000",
31753 => "0000000000000000",31754 => "0000000000000000",
31755 => "0000000000000000",31756 => "0000000000000000",
31757 => "0000000000000000",31758 => "0000000000000000",
31759 => "0000000000000000",31760 => "0000000000000000",
31761 => "0000000000000000",31762 => "0000000000000000",
31763 => "0000000000000000",31764 => "0000000000000000",
31765 => "0000000000000000",31766 => "0000000000000000",
31767 => "0000000000000000",31768 => "0000000000000000",
31769 => "0000000000000000",31770 => "0000000000000000",
31771 => "0000000000000000",31772 => "0000000000000000",
31773 => "0000000000000000",31774 => "0000000000000000",
31775 => "0000000000000000",31776 => "0000000000000000",
31777 => "0000000000000000",31778 => "0000000000000000",
31779 => "0000000000000000",31780 => "0000000000000000",
31781 => "0000000000000000",31782 => "0000000000000000",
31783 => "0000000000000000",31784 => "0000000000000000",
31785 => "0000000000000000",31786 => "0000000000000000",
31787 => "0000000000000000",31788 => "0000000000000000",
31789 => "0000000000000000",31790 => "0000000000000000",
31791 => "0000000000000000",31792 => "0000000000000000",
31793 => "0000000000000000",31794 => "0000000000000000",
31795 => "0000000000000000",31796 => "0000000000000000",
31797 => "0000000000000000",31798 => "0000000000000000",
31799 => "0000000000000000",31800 => "0000000000000000",
31801 => "0000000000000000",31802 => "0000000000000000",
31803 => "0000000000000000",31804 => "0000000000000000",
31805 => "0000000000000000",31806 => "0000000000000000",
31807 => "0000000000000000",31808 => "0000000000000000",
31809 => "0000000000000000",31810 => "0000000000000000",
31811 => "0000000000000000",31812 => "0000000000000000",
31813 => "0000000000000000",31814 => "0000000000000000",
31815 => "0000000000000000",31816 => "0000000000000000",
31817 => "0000000000000000",31818 => "0000000000000000",
31819 => "0000000000000000",31820 => "0000000000000000",
31821 => "0000000000000000",31822 => "0000000000000000",
31823 => "0000000000000000",31824 => "0000000000000000",
31825 => "0000000000000000",31826 => "0000000000000000",
31827 => "0000000000000000",31828 => "0000000000000000",
31829 => "0000000000000000",31830 => "0000000000000000",
31831 => "0000000000000000",31832 => "0000000000000000",
31833 => "0000000000000000",31834 => "0000000000000000",
31835 => "0000000000000000",31836 => "0000000000000000",
31837 => "0000000000000000",31838 => "0000000000000000",
31839 => "0000000000000000",31840 => "0000000000000000",
31841 => "0000000000000000",31842 => "0000000000000000",
31843 => "0000000000000000",31844 => "0000000000000000",
31845 => "0000000000000000",31846 => "0000000000000000",
31847 => "0000000000000000",31848 => "0000000000000000",
31849 => "0000000000000000",31850 => "0000000000000000",
31851 => "0000000000000000",31852 => "0000000000000000",
31853 => "0000000000000000",31854 => "0000000000000000",
31855 => "0000000000000000",31856 => "0000000000000000",
31857 => "0000000000000000",31858 => "0000000000000000",
31859 => "0000000000000000",31860 => "0000000000000000",
31861 => "0000000000000000",31862 => "0000000000000000",
31863 => "0000000000000000",31864 => "0000000000000000",
31865 => "0000000000000000",31866 => "0000000000000000",
31867 => "0000000000000000",31868 => "0000000000000000",
31869 => "0000000000000000",31870 => "0000000000000000",
31871 => "0000000000000000",31872 => "0000000000000000",
31873 => "0000000000000000",31874 => "0000000000000000",
31875 => "0000000000000000",31876 => "0000000000000000",
31877 => "0000000000000000",31878 => "0000000000000000",
31879 => "0000000000000000",31880 => "0000000000000000",
31881 => "0000000000000000",31882 => "0000000000000000",
31883 => "0000000000000000",31884 => "0000000000000000",
31885 => "0000000000000000",31886 => "0000000000000000",
31887 => "0000000000000000",31888 => "0000000000000000",
31889 => "0000000000000000",31890 => "0000000000000000",
31891 => "0000000000000000",31892 => "0000000000000000",
31893 => "0000000000000000",31894 => "0000000000000000",
31895 => "0000000000000000",31896 => "0000000000000000",
31897 => "0000000000000000",31898 => "0000000000000000",
31899 => "0000000000000000",31900 => "0000000000000000",
31901 => "0000000000000000",31902 => "0000000000000000",
31903 => "0000000000000000",31904 => "0000000000000000",
31905 => "0000000000000000",31906 => "0000000000000000",
31907 => "0000000000000000",31908 => "0000000000000000",
31909 => "0000000000000000",31910 => "0000000000000000",
31911 => "0000000000000000",31912 => "0000000000000000",
31913 => "0000000000000000",31914 => "0000000000000000",
31915 => "0000000000000000",31916 => "0000000000000000",
31917 => "0000000000000000",31918 => "0000000000000000",
31919 => "0000000000000000",31920 => "0000000000000000",
31921 => "0000000000000000",31922 => "0000000000000000",
31923 => "0000000000000000",31924 => "0000000000000000",
31925 => "0000000000000000",31926 => "0000000000000000",
31927 => "0000000000000000",31928 => "0000000000000000",
31929 => "0000000000000000",31930 => "0000000000000000",
31931 => "0000000000000000",31932 => "0000000000000000",
31933 => "0000000000000000",31934 => "0000000000000000",
31935 => "0000000000000000",31936 => "0000000000000000",
31937 => "0000000000000000",31938 => "0000000000000000",
31939 => "0000000000000000",31940 => "0000000000000000",
31941 => "0000000000000000",31942 => "0000000000000000",
31943 => "0000000000000000",31944 => "0000000000000000",
31945 => "0000000000000000",31946 => "0000000000000000",
31947 => "0000000000000000",31948 => "0000000000000000",
31949 => "0000000000000000",31950 => "0000000000000000",
31951 => "0000000000000000",31952 => "0000000000000000",
31953 => "0000000000000000",31954 => "0000000000000000",
31955 => "0000000000000000",31956 => "0000000000000000",
31957 => "0000000000000000",31958 => "0000000000000000",
31959 => "0000000000000000",31960 => "0000000000000000",
31961 => "0000000000000000",31962 => "0000000000000000",
31963 => "0000000000000000",31964 => "0000000000000000",
31965 => "0000000000000000",31966 => "0000000000000000",
31967 => "0000000000000000",31968 => "0000000000000000",
31969 => "0000000000000000",31970 => "0000000000000000",
31971 => "0000000000000000",31972 => "0000000000000000",
31973 => "0000000000000000",31974 => "0000000000000000",
31975 => "0000000000000000",31976 => "0000000000000000",
31977 => "0000000000000000",31978 => "0000000000000000",
31979 => "0000000000000000",31980 => "0000000000000000",
31981 => "0000000000000000",31982 => "0000000000000000",
31983 => "0000000000000000",31984 => "0000000000000000",
31985 => "0000000000000000",31986 => "0000000000000000",
31987 => "0000000000000000",31988 => "0000000000000000",
31989 => "0000000000000000",31990 => "0000000000000000",
31991 => "0000000000000000",31992 => "0000000000000000",
31993 => "0000000000000000",31994 => "0000000000000000",
31995 => "0000000000000000",31996 => "0000000000000000",
31997 => "0000000000000000",31998 => "0000000000000000",
31999 => "0000000000000000",32000 => "0000000000000000",
32001 => "0000000000000000",32002 => "0000000000000000",
32003 => "0000000000000000",32004 => "0000000000000000",
32005 => "0000000000000000",32006 => "0000000000000000",
32007 => "0000000000000000",32008 => "0000000000000000",
32009 => "0000000000000000",32010 => "0000000000000000",
32011 => "0000000000000000",32012 => "0000000000000000",
32013 => "0000000000000000",32014 => "0000000000000000",
32015 => "0000000000000000",32016 => "0000000000000000",
32017 => "0000000000000000",32018 => "0000000000000000",
32019 => "0000000000000000",32020 => "0000000000000000",
32021 => "0000000000000000",32022 => "0000000000000000",
32023 => "0000000000000000",32024 => "0000000000000000",
32025 => "0000000000000000",32026 => "0000000000000000",
32027 => "0000000000000000",32028 => "0000000000000000",
32029 => "0000000000000000",32030 => "0000000000000000",
32031 => "0000000000000000",32032 => "0000000000000000",
32033 => "0000000000000000",32034 => "0000000000000000",
32035 => "0000000000000000",32036 => "0000000000000000",
32037 => "0000000000000000",32038 => "0000000000000000",
32039 => "0000000000000000",32040 => "0000000000000000",
32041 => "0000000000000000",32042 => "0000000000000000",
32043 => "0000000000000000",32044 => "0000000000000000",
32045 => "0000000000000000",32046 => "0000000000000000",
32047 => "0000000000000000",32048 => "0000000000000000",
32049 => "0000000000000000",32050 => "0000000000000000",
32051 => "0000000000000000",32052 => "0000000000000000",
32053 => "0000000000000000",32054 => "0000000000000000",
32055 => "0000000000000000",32056 => "0000000000000000",
32057 => "0000000000000000",32058 => "0000000000000000",
32059 => "0000000000000000",32060 => "0000000000000000",
32061 => "0000000000000000",32062 => "0000000000000000",
32063 => "0000000000000000",32064 => "0000000000000000",
32065 => "0000000000000000",32066 => "0000000000000000",
32067 => "0000000000000000",32068 => "0000000000000000",
32069 => "0000000000000000",32070 => "0000000000000000",
32071 => "0000000000000000",32072 => "0000000000000000",
32073 => "0000000000000000",32074 => "0000000000000000",
32075 => "0000000000000000",32076 => "0000000000000000",
32077 => "0000000000000000",32078 => "0000000000000000",
32079 => "0000000000000000",32080 => "0000000000000000",
32081 => "0000000000000000",32082 => "0000000000000000",
32083 => "0000000000000000",32084 => "0000000000000000",
32085 => "0000000000000000",32086 => "0000000000000000",
32087 => "0000000000000000",32088 => "0000000000000000",
32089 => "0000000000000000",32090 => "0000000000000000",
32091 => "0000000000000000",32092 => "0000000000000000",
32093 => "0000000000000000",32094 => "0000000000000000",
32095 => "0000000000000000",32096 => "0000000000000000",
32097 => "0000000000000000",32098 => "0000000000000000",
32099 => "0000000000000000",32100 => "0000000000000000",
32101 => "0000000000000000",32102 => "0000000000000000",
32103 => "0000000000000000",32104 => "0000000000000000",
32105 => "0000000000000000",32106 => "0000000000000000",
32107 => "0000000000000000",32108 => "0000000000000000",
32109 => "0000000000000000",32110 => "0000000000000000",
32111 => "0000000000000000",32112 => "0000000000000000",
32113 => "0000000000000000",32114 => "0000000000000000",
32115 => "0000000000000000",32116 => "0000000000000000",
32117 => "0000000000000000",32118 => "0000000000000000",
32119 => "0000000000000000",32120 => "0000000000000000",
32121 => "0000000000000000",32122 => "0000000000000000",
32123 => "0000000000000000",32124 => "0000000000000000",
32125 => "0000000000000000",32126 => "0000000000000000",
32127 => "0000000000000000",32128 => "0000000000000000",
32129 => "0000000000000000",32130 => "0000000000000000",
32131 => "0000000000000000",32132 => "0000000000000000",
32133 => "0000000000000000",32134 => "0000000000000000",
32135 => "0000000000000000",32136 => "0000000000000000",
32137 => "0000000000000000",32138 => "0000000000000000",
32139 => "0000000000000000",32140 => "0000000000000000",
32141 => "0000000000000000",32142 => "0000000000000000",
32143 => "0000000000000000",32144 => "0000000000000000",
32145 => "0000000000000000",32146 => "0000000000000000",
32147 => "0000000000000000",32148 => "0000000000000000",
32149 => "0000000000000000",32150 => "0000000000000000",
32151 => "0000000000000000",32152 => "0000000000000000",
32153 => "0000000000000000",32154 => "0000000000000000",
32155 => "0000000000000000",32156 => "0000000000000000",
32157 => "0000000000000000",32158 => "0000000000000000",
32159 => "0000000000000000",32160 => "0000000000000000",
32161 => "0000000000000000",32162 => "0000000000000000",
32163 => "0000000000000000",32164 => "0000000000000000",
32165 => "0000000000000000",32166 => "0000000000000000",
32167 => "0000000000000000",32168 => "0000000000000000",
32169 => "0000000000000000",32170 => "0000000000000000",
32171 => "0000000000000000",32172 => "0000000000000000",
32173 => "0000000000000000",32174 => "0000000000000000",
32175 => "0000000000000000",32176 => "0000000000000000",
32177 => "0000000000000000",32178 => "0000000000000000",
32179 => "0000000000000000",32180 => "0000000000000000",
32181 => "0000000000000000",32182 => "0000000000000000",
32183 => "0000000000000000",32184 => "0000000000000000",
32185 => "0000000000000000",32186 => "0000000000000000",
32187 => "0000000000000000",32188 => "0000000000000000",
32189 => "0000000000000000",32190 => "0000000000000000",
32191 => "0000000000000000",32192 => "0000000000000000",
32193 => "0000000000000000",32194 => "0000000000000000",
32195 => "0000000000000000",32196 => "0000000000000000",
32197 => "0000000000000000",32198 => "0000000000000000",
32199 => "0000000000000000",32200 => "0000000000000000",
32201 => "0000000000000000",32202 => "0000000000000000",
32203 => "0000000000000000",32204 => "0000000000000000",
32205 => "0000000000000000",32206 => "0000000000000000",
32207 => "0000000000000000",32208 => "0000000000000000",
32209 => "0000000000000000",32210 => "0000000000000000",
32211 => "0000000000000000",32212 => "0000000000000000",
32213 => "0000000000000000",32214 => "0000000000000000",
32215 => "0000000000000000",32216 => "0000000000000000",
32217 => "0000000000000000",32218 => "0000000000000000",
32219 => "0000000000000000",32220 => "0000000000000000",
32221 => "0000000000000000",32222 => "0000000000000000",
32223 => "0000000000000000",32224 => "0000000000000000",
32225 => "0000000000000000",32226 => "0000000000000000",
32227 => "0000000000000000",32228 => "0000000000000000",
32229 => "0000000000000000",32230 => "0000000000000000",
32231 => "0000000000000000",32232 => "0000000000000000",
32233 => "0000000000000000",32234 => "0000000000000000",
32235 => "0000000000000000",32236 => "0000000000000000",
32237 => "0000000000000000",32238 => "0000000000000000",
32239 => "0000000000000000",32240 => "0000000000000000",
32241 => "0000000000000000",32242 => "0000000000000000",
32243 => "0000000000000000",32244 => "0000000000000000",
32245 => "0000000000000000",32246 => "0000000000000000",
32247 => "0000000000000000",32248 => "0000000000000000",
32249 => "0000000000000000",32250 => "0000000000000000",
32251 => "0000000000000000",32252 => "0000000000000000",
32253 => "0000000000000000",32254 => "0000000000000000",
32255 => "0000000000000000",32256 => "0000000000000000",
32257 => "0000000000000000",32258 => "0000000000000000",
32259 => "0000000000000000",32260 => "0000000000000000",
32261 => "0000000000000000",32262 => "0000000000000000",
32263 => "0000000000000000",32264 => "0000000000000000",
32265 => "0000000000000000",32266 => "0000000000000000",
32267 => "0000000000000000",32268 => "0000000000000000",
32269 => "0000000000000000",32270 => "0000000000000000",
32271 => "0000000000000000",32272 => "0000000000000000",
32273 => "0000000000000000",32274 => "0000000000000000",
32275 => "0000000000000000",32276 => "0000000000000000",
32277 => "0000000000000000",32278 => "0000000000000000",
32279 => "0000000000000000",32280 => "0000000000000000",
32281 => "0000000000000000",32282 => "0000000000000000",
32283 => "0000000000000000",32284 => "0000000000000000",
32285 => "0000000000000000",32286 => "0000000000000000",
32287 => "0000000000000000",32288 => "0000000000000000",
32289 => "0000000000000000",32290 => "0000000000000000",
32291 => "0000000000000000",32292 => "0000000000000000",
32293 => "0000000000000000",32294 => "0000000000000000",
32295 => "0000000000000000",32296 => "0000000000000000",
32297 => "0000000000000000",32298 => "0000000000000000",
32299 => "0000000000000000",32300 => "0000000000000000",
32301 => "0000000000000000",32302 => "0000000000000000",
32303 => "0000000000000000",32304 => "0000000000000000",
32305 => "0000000000000000",32306 => "0000000000000000",
32307 => "0000000000000000",32308 => "0000000000000000",
32309 => "0000000000000000",32310 => "0000000000000000",
32311 => "0000000000000000",32312 => "0000000000000000",
32313 => "0000000000000000",32314 => "0000000000000000",
32315 => "0000000000000000",32316 => "0000000000000000",
32317 => "0000000000000000",32318 => "0000000000000000",
32319 => "0000000000000000",32320 => "0000000000000000",
32321 => "0000000000000000",32322 => "0000000000000000",
32323 => "0000000000000000",32324 => "0000000000000000",
32325 => "0000000000000000",32326 => "0000000000000000",
32327 => "0000000000000000",32328 => "0000000000000000",
32329 => "0000000000000000",32330 => "0000000000000000",
32331 => "0000000000000000",32332 => "0000000000000000",
32333 => "0000000000000000",32334 => "0000000000000000",
32335 => "0000000000000000",32336 => "0000000000000000",
32337 => "0000000000000000",32338 => "0000000000000000",
32339 => "0000000000000000",32340 => "0000000000000000",
32341 => "0000000000000000",32342 => "0000000000000000",
32343 => "0000000000000000",32344 => "0000000000000000",
32345 => "0000000000000000",32346 => "0000000000000000",
32347 => "0000000000000000",32348 => "0000000000000000",
32349 => "0000000000000000",32350 => "0000000000000000",
32351 => "0000000000000000",32352 => "0000000000000000",
32353 => "0000000000000000",32354 => "0000000000000000",
32355 => "0000000000000000",32356 => "0000000000000000",
32357 => "0000000000000000",32358 => "0000000000000000",
32359 => "0000000000000000",32360 => "0000000000000000",
32361 => "0000000000000000",32362 => "0000000000000000",
32363 => "0000000000000000",32364 => "0000000000000000",
32365 => "0000000000000000",32366 => "0000000000000000",
32367 => "0000000000000000",32368 => "0000000000000000",
32369 => "0000000000000000",32370 => "0000000000000000",
32371 => "0000000000000000",32372 => "0000000000000000",
32373 => "0000000000000000",32374 => "0000000000000000",
32375 => "0000000000000000",32376 => "0000000000000000",
32377 => "0000000000000000",32378 => "0000000000000000",
32379 => "0000000000000000",32380 => "0000000000000000",
32381 => "0000000000000000",32382 => "0000000000000000",
32383 => "0000000000000000",32384 => "0000000000000000",
32385 => "0000000000000000",32386 => "0000000000000000",
32387 => "0000000000000000",32388 => "0000000000000000",
32389 => "0000000000000000",32390 => "0000000000000000",
32391 => "0000000000000000",32392 => "0000000000000000",
32393 => "0000000000000000",32394 => "0000000000000000",
32395 => "0000000000000000",32396 => "0000000000000000",
32397 => "0000000000000000",32398 => "0000000000000000",
32399 => "0000000000000000",32400 => "0000000000000000",
32401 => "0000000000000000",32402 => "0000000000000000",
32403 => "0000000000000000",32404 => "0000000000000000",
32405 => "0000000000000000",32406 => "0000000000000000",
32407 => "0000000000000000",32408 => "0000000000000000",
32409 => "0000000000000000",32410 => "0000000000000000",
32411 => "0000000000000000",32412 => "0000000000000000",
32413 => "0000000000000000",32414 => "0000000000000000",
32415 => "0000000000000000",32416 => "0000000000000000",
32417 => "0000000000000000",32418 => "0000000000000000",
32419 => "0000000000000000",32420 => "0000000000000000",
32421 => "0000000000000000",32422 => "0000000000000000",
32423 => "0000000000000000",32424 => "0000000000000000",
32425 => "0000000000000000",32426 => "0000000000000000",
32427 => "0000000000000000",32428 => "0000000000000000",
32429 => "0000000000000000",32430 => "0000000000000000",
32431 => "0000000000000000",32432 => "0000000000000000",
32433 => "0000000000000000",32434 => "0000000000000000",
32435 => "0000000000000000",32436 => "0000000000000000",
32437 => "0000000000000000",32438 => "0000000000000000",
32439 => "0000000000000000",32440 => "0000000000000000",
32441 => "0000000000000000",32442 => "0000000000000000",
32443 => "0000000000000000",32444 => "0000000000000000",
32445 => "0000000000000000",32446 => "0000000000000000",
32447 => "0000000000000000",32448 => "0000000000000000",
32449 => "0000000000000000",32450 => "0000000000000000",
32451 => "0000000000000000",32452 => "0000000000000000",
32453 => "0000000000000000",32454 => "0000000000000000",
32455 => "0000000000000000",32456 => "0000000000000000",
32457 => "0000000000000000",32458 => "0000000000000000",
32459 => "0000000000000000",32460 => "0000000000000000",
32461 => "0000000000000000",32462 => "0000000000000000",
32463 => "0000000000000000",32464 => "0000000000000000",
32465 => "0000000000000000",32466 => "0000000000000000",
32467 => "0000000000000000",32468 => "0000000000000000",
32469 => "0000000000000000",32470 => "0000000000000000",
32471 => "0000000000000000",32472 => "0000000000000000",
32473 => "0000000000000000",32474 => "0000000000000000",
32475 => "0000000000000000",32476 => "0000000000000000",
32477 => "0000000000000000",32478 => "0000000000000000",
32479 => "0000000000000000",32480 => "0000000000000000",
32481 => "0000000000000000",32482 => "0000000000000000",
32483 => "0000000000000000",32484 => "0000000000000000",
32485 => "0000000000000000",32486 => "0000000000000000",
32487 => "0000000000000000",32488 => "0000000000000000",
32489 => "0000000000000000",32490 => "0000000000000000",
32491 => "0000000000000000",32492 => "0000000000000000",
32493 => "0000000000000000",32494 => "0000000000000000",
32495 => "0000000000000000",32496 => "0000000000000000",
32497 => "0000000000000000",32498 => "0000000000000000",
32499 => "0000000000000000",32500 => "0000000000000000",
32501 => "0000000000000000",32502 => "0000000000000000",
32503 => "0000000000000000",32504 => "0000000000000000",
32505 => "0000000000000000",32506 => "0000000000000000",
32507 => "0000000000000000",32508 => "0000000000000000",
32509 => "0000000000000000",32510 => "0000000000000000",
32511 => "0000000000000000",32512 => "0000000000000000",
32513 => "0000000000000000",32514 => "0000000000000000",
32515 => "0000000000000000",32516 => "0000000000000000",
32517 => "0000000000000000",32518 => "0000000000000000",
32519 => "0000000000000000",32520 => "0000000000000000",
32521 => "0000000000000000",32522 => "0000000000000000",
32523 => "0000000000000000",32524 => "0000000000000000",
32525 => "0000000000000000",32526 => "0000000000000000",
32527 => "0000000000000000",32528 => "0000000000000000",
32529 => "0000000000000000",32530 => "0000000000000000",
32531 => "0000000000000000",32532 => "0000000000000000",
32533 => "0000000000000000",32534 => "0000000000000000",
32535 => "0000000000000000",32536 => "0000000000000000",
32537 => "0000000000000000",32538 => "0000000000000000",
32539 => "0000000000000000",32540 => "0000000000000000",
32541 => "0000000000000000",32542 => "0000000000000000",
32543 => "0000000000000000",32544 => "0000000000000000",
32545 => "0000000000000000",32546 => "0000000000000000",
32547 => "0000000000000000",32548 => "0000000000000000",
32549 => "0000000000000000",32550 => "0000000000000000",
32551 => "0000000000000000",32552 => "0000000000000000",
32553 => "0000000000000000",32554 => "0000000000000000",
32555 => "0000000000000000",32556 => "0000000000000000",
32557 => "0000000000000000",32558 => "0000000000000000",
32559 => "0000000000000000",32560 => "0000000000000000",
32561 => "0000000000000000",32562 => "0000000000000000",
32563 => "0000000000000000",32564 => "0000000000000000",
32565 => "0000000000000000",32566 => "0000000000000000",
32567 => "0000000000000000",32568 => "0000000000000000",
32569 => "0000000000000000",32570 => "0000000000000000",
32571 => "0000000000000000",32572 => "0000000000000000",
32573 => "0000000000000000",32574 => "0000000000000000",
32575 => "0000000000000000",32576 => "0000000000000000",
32577 => "0000000000000000",32578 => "0000000000000000",
32579 => "0000000000000000",32580 => "0000000000000000",
32581 => "0000000000000000",32582 => "0000000000000000",
32583 => "0000000000000000",32584 => "0000000000000000",
32585 => "0000000000000000",32586 => "0000000000000000",
32587 => "0000000000000000",32588 => "0000000000000000",
32589 => "0000000000000000",32590 => "0000000000000000",
32591 => "0000000000000000",32592 => "0000000000000000",
32593 => "0000000000000000",32594 => "0000000000000000",
32595 => "0000000000000000",32596 => "0000000000000000",
32597 => "0000000000000000",32598 => "0000000000000000",
32599 => "0000000000000000",32600 => "0000000000000000",
32601 => "0000000000000000",32602 => "0000000000000000",
32603 => "0000000000000000",32604 => "0000000000000000",
32605 => "0000000000000000",32606 => "0000000000000000",
32607 => "0000000000000000",32608 => "0000000000000000",
32609 => "0000000000000000",32610 => "0000000000000000",
32611 => "0000000000000000",32612 => "0000000000000000",
32613 => "0000000000000000",32614 => "0000000000000000",
32615 => "0000000000000000",32616 => "0000000000000000",
32617 => "0000000000000000",32618 => "0000000000000000",
32619 => "0000000000000000",32620 => "0000000000000000",
32621 => "0000000000000000",32622 => "0000000000000000",
32623 => "0000000000000000",32624 => "0000000000000000",
32625 => "0000000000000000",32626 => "0000000000000000",
32627 => "0000000000000000",32628 => "0000000000000000",
32629 => "0000000000000000",32630 => "0000000000000000",
32631 => "0000000000000000",32632 => "0000000000000000",
32633 => "0000000000000000",32634 => "0000000000000000",
32635 => "0000000000000000",32636 => "0000000000000000",
32637 => "0000000000000000",32638 => "0000000000000000",
32639 => "0000000000000000",32640 => "0000000000000000",
32641 => "0000000000000000",32642 => "0000000000000000",
32643 => "0000000000000000",32644 => "0000000000000000",
32645 => "0000000000000000",32646 => "0000000000000000",
32647 => "0000000000000000",32648 => "0000000000000000",
32649 => "0000000000000000",32650 => "0000000000000000",
32651 => "0000000000000000",32652 => "0000000000000000",
32653 => "0000000000000000",32654 => "0000000000000000",
32655 => "0000000000000000",32656 => "0000000000000000",
32657 => "0000000000000000",32658 => "0000000000000000",
32659 => "0000000000000000",32660 => "0000000000000000",
32661 => "0000000000000000",32662 => "0000000000000000",
32663 => "0000000000000000",32664 => "0000000000000000",
32665 => "0000000000000000",32666 => "0000000000000000",
32667 => "0000000000000000",32668 => "0000000000000000",
32669 => "0000000000000000",32670 => "0000000000000000",
32671 => "0000000000000000",32672 => "0000000000000000",
32673 => "0000000000000000",32674 => "0000000000000000",
32675 => "0000000000000000",32676 => "0000000000000000",
32677 => "0000000000000000",32678 => "0000000000000000",
32679 => "0000000000000000",32680 => "0000000000000000",
32681 => "0000000000000000",32682 => "0000000000000000",
32683 => "0000000000000000",32684 => "0000000000000000",
32685 => "0000000000000000",32686 => "0000000000000000",
32687 => "0000000000000000",32688 => "0000000000000000",
32689 => "0000000000000000",32690 => "0000000000000000",
32691 => "0000000000000000",32692 => "0000000000000000",
32693 => "0000000000000000",32694 => "0000000000000000",
32695 => "0000000000000000",32696 => "0000000000000000",
32697 => "0000000000000000",32698 => "0000000000000000",
32699 => "0000000000000000",32700 => "0000000000000000",
32701 => "0000000000000000",32702 => "0000000000000000",
32703 => "0000000000000000",32704 => "0000000000000000",
32705 => "0000000000000000",32706 => "0000000000000000",
32707 => "0000000000000000",32708 => "0000000000000000",
32709 => "0000000000000000",32710 => "0000000000000000",
32711 => "0000000000000000",32712 => "0000000000000000",
32713 => "0000000000000000",32714 => "0000000000000000",
32715 => "0000000000000000",32716 => "0000000000000000",
32717 => "0000000000000000",32718 => "0000000000000000",
32719 => "0000000000000000",32720 => "0000000000000000",
32721 => "0000000000000000",32722 => "0000000000000000",
32723 => "0000000000000000",32724 => "0000000000000000",
32725 => "0000000000000000",32726 => "0000000000000000",
32727 => "0000000000000000",32728 => "0000000000000000",
32729 => "0000000000000000",32730 => "0000000000000000",
32731 => "0000000000000000",32732 => "0000000000000000",
32733 => "0000000000000000",32734 => "0000000000000000",
32735 => "0000000000000000",32736 => "0000000000000000",
32737 => "0000000000000000",32738 => "0000000000000000",
32739 => "0000000000000000",32740 => "0000000000000000",
32741 => "0000000000000000",32742 => "0000000000000000",
32743 => "0000000000000000",32744 => "0000000000000000",
32745 => "0000000000000000",32746 => "0000000000000000",
32747 => "0000000000000000",32748 => "0000000000000000",
32749 => "0000000000000000",32750 => "0000000000000000",
32751 => "0000000000000000",32752 => "0000000000000000",
32753 => "0000000000000000",32754 => "0000000000000000",
32755 => "0000000000000000",32756 => "0000000000000000",
32757 => "0000000000000000",32758 => "0000000000000000",
32759 => "0000000000000000",32760 => "0000000000000000",
32761 => "0000000000000000",32762 => "0000000000000000",
32763 => "0000000000000000",32764 => "0000000000000000",
32765 => "0000000000000000",32766 => "0000000000000000",
32767 => "0000000000000000",32768 => "0000100000000000",
32769 => "0000001110001001",32770 => "0000001100110011",
32771 => "0000001011100101",32772 => "0000000001000011",
32773 => "0000001001011111",32774 => "0000001000100101",
32775 => "0000000111110001",32776 => "0000000111000001",
32777 => "0000000110010111",32778 => "0000001110001001",
32779 => "0000001110000000",32780 => "0000001101110111",
32781 => "0000001101101110",32782 => "0000001101100101",
32783 => "0000001101011101",32784 => "0000001101010100",
32785 => "0000001101001100",32786 => "0000001101000011",
32787 => "0000001100111011",32788 => "0000001100110011",
32789 => "0000001100101011",32790 => "0000001100100011",
32791 => "0000001100011011",32792 => "0000001100010011",
32793 => "0000001100001011",32794 => "0000001100000011",
32795 => "0000001011111011",32796 => "0000001011110100",
32797 => "0000001011101100",32798 => "0000001011100101",
32799 => "0000001011011101",32800 => "0000001011010110",
32801 => "0000001011001111",32802 => "0000001011001000",
32803 => "0000001011000001",32804 => "0000001010111010",
32805 => "0000001010110011",32806 => "0000001010101100",
32807 => "0000001010100101",32808 => "0000000001000011",
32809 => "0000001010011000",32810 => "0000001010010001",
32811 => "0000001010001011",32812 => "0000001010000100",
32813 => "0000001001111110",32814 => "0000001001110111",
32815 => "0000001001110001",32816 => "0000001001101011",
32817 => "0000001001100101",32818 => "0000001001011111",
32819 => "0000000000000110",32820 => "0000001001010011",
32821 => "0000001001001101",32822 => "0000001001000111",
32823 => "0000001001000001",32824 => "0000001000111011",
32825 => "0000001000110110",32826 => "0000000000111000",
32827 => "0000001000101010",32828 => "0000001000100101",
32829 => "0000001000011111",32830 => "0000001000011010",
32831 => "0000001000010101",32832 => "0000001000001111",
32833 => "0000001000001010",32834 => "0000001000000101",
32835 => "0000001000000000",32836 => "0000000111111011",
32837 => "0000000111110110",32838 => "0000000111110001",
32839 => "0000000111101100",32840 => "0000000111100111",
32841 => "0000000111100010",32842 => "0000000111011101",
32843 => "0000000111011000",32844 => "0000000111010100",
32845 => "0000000111001111",32846 => "0000000111001010",
32847 => "0000000111000110",32848 => "0000000111000001",
32849 => "0000000110111101",32850 => "0000000000101100",
32851 => "0000000110110100",32852 => "0000000110110000",
32853 => "0000000110101011",32854 => "0000000110100111",
32855 => "0000000110100011",32856 => "0000000110011111",
32857 => "0000000110011011",32858 => "0000000110010111",
32859 => "0000000110010011",32860 => "0000000110001111",
32861 => "0000000110001011",32862 => "0000000110000111",
32863 => "0000000110000011",32864 => "0000000101111111",
32865 => "0000000101111011",32866 => "0000000101110111",
32867 => "0000000101110100",32868 => "0000001110001001",
32869 => "0000001110001000",32870 => "0000001110000111",
32871 => "0000001110000110",32872 => "0000001110000101",
32873 => "0000000000001001",32874 => "0000001110000011",
32875 => "0000001110000011",32876 => "0000001110000010",
32877 => "0000001110000001",32878 => "0000001110000000",
32879 => "0000001101111111",32880 => "0000001101111110",
32881 => "0000001101111101",32882 => "0000001101111100",
32883 => "0000001101111011",32884 => "0000000001011001",
32885 => "0000000001011001",32886 => "0000001101111001",
32887 => "0000001101111000",32888 => "0000001101110111",
32889 => "0000001101110110",32890 => "0000001101110101",
32891 => "0000001101110100",32892 => "0000001101110011",
32893 => "0000001101110010",32894 => "0000001101110010",
32895 => "0000001101110001",32896 => "0000000001011000",
32897 => "0000001101101111",32898 => "0000001101101110",
32899 => "0000001101101101",32900 => "0000001101101100",
32901 => "0000001101101011",32902 => "0000001101101011",
32903 => "0000001101101010",32904 => "0000001101101001",
32905 => "0000001101101000",32906 => "0000001101100111",
32907 => "0000000001010111",32908 => "0000001101100101",
32909 => "0000001101100100",32910 => "0000001101100100",
32911 => "0000001101100011",32912 => "0000001101100010",
32913 => "0000001101100001",32914 => "0000001101100000",
32915 => "0000001101011111",32916 => "0000001101011110",
32917 => "0000001101011110",32918 => "0000001101011101",
32919 => "0000000001010110",32920 => "0000001101011011",
32921 => "0000001101011010",32922 => "0000001101011001",
32923 => "0000001101011000",32924 => "0000001101011000",
32925 => "0000001101010111",32926 => "0000001101010110",
32927 => "0000001101010101",32928 => "0000001101010100",
32929 => "0000001101010011",32930 => "0000000001010101",
32931 => "0000000001010101",32932 => "0000001101010001",
32933 => "0000001101010000",32934 => "0000001101001111",
32935 => "0000001101001110",32936 => "0000001101001101",
32937 => "0000001101001101",32938 => "0000001101001100",
32939 => "0000001101001011",32940 => "0000001101001010",
32941 => "0000001101001001",32942 => "0000000001010100",
32943 => "0000001101000111",32944 => "0000001101000111",
32945 => "0000001101000110",32946 => "0000001101000101",
32947 => "0000001101000100",32948 => "0000001101000011",
32949 => "0000001101000010",32950 => "0000001101000010",
32951 => "0000001101000001",32952 => "0000001101000000",
32953 => "0000001100111111",32954 => "0000000001010011",
32955 => "0000001100111101",32956 => "0000001100111101",
32957 => "0000001100111100",32958 => "0000001100111011",
32959 => "0000001100111010",32960 => "0000001100111001",
32961 => "0000001100111000",32962 => "0000001100111000",
32963 => "0000001100110111",32964 => "0000001100110110",
32965 => "0000001100110101",32966 => "0000000001010010",
32967 => "0000000001010010",32968 => "0000001100110011",
32969 => "0000001100110010",32970 => "0000001100110001",
32971 => "0000001100110000",32972 => "0000001100101111",
32973 => "0000001100101111",32974 => "0000001100101110",
32975 => "0000001100101101",32976 => "0000001100101100",
32977 => "0000001100101011",32978 => "0000001100101011",
32979 => "0000000001010001",32980 => "0000001100101001",
32981 => "0000001100101000",32982 => "0000001100100111",
32983 => "0000001100100111",32984 => "0000001100100110",
32985 => "0000001100100101",32986 => "0000001100100100",
32987 => "0000001100100011",32988 => "0000001100100011",
32989 => "0000001100100010",32990 => "0000001100100001",
32991 => "0000000000001000",32992 => "0000001100011111",
32993 => "0000001100011111",32994 => "0000001100011110",
32995 => "0000001100011101",32996 => "0000001100011100",
32997 => "0000001100011011",32998 => "0000001100011011",
32999 => "0000001100011010",33000 => "0000001100011001",
33001 => "0000001100011000",33002 => "0000001100010111",
33003 => "0000001100010111",33004 => "0000000001001111",
33005 => "0000001100010101",33006 => "0000001100010100",
33007 => "0000001100010011",33008 => "0000001100010011",
33009 => "0000001100010010",33010 => "0000001100010001",
33011 => "0000001100010000",33012 => "0000001100001111",
33013 => "0000001100001111",33014 => "0000001100001110",
33015 => "0000001100001101",33016 => "0000000001001110",
33017 => "0000000001001110",33018 => "0000001100001011",
33019 => "0000001100001010",33020 => "0000001100001001",
33021 => "0000001100001000",33022 => "0000001100001000",
33023 => "0000001100000111",33024 => "0000001100000110",
33025 => "0000001100000101",33026 => "0000001100000101",
33027 => "0000001100000100",33028 => "0000001100000011",
33029 => "0000000001001101",33030 => "0000000001001101",
33031 => "0000001100000001",33032 => "0000001100000000",
33033 => "0000001011111111",33034 => "0000001011111110",
33035 => "0000001011111110",33036 => "0000001011111101",
33037 => "0000001011111100",33038 => "0000001011111011",
33039 => "0000001011111011",33040 => "0000001011111010",
33041 => "0000001011111001",33042 => "0000000001001100",
33043 => "0000000001001100",33044 => "0000001011110111",
33045 => "0000001011110110",33046 => "0000001011110101",
33047 => "0000001011110101",33048 => "0000001011110100",
33049 => "0000001011110011",33050 => "0000001011110010",
33051 => "0000001011110010",33052 => "0000001011110001",
33053 => "0000001011110000",33054 => "0000001011101111",
33055 => "0000001011101111",33056 => "0000000001001011",
33057 => "0000001011101101",33058 => "0000001011101100",
33059 => "0000001011101100",33060 => "0000001011101011",
33061 => "0000001011101010",33062 => "0000001011101001",
33063 => "0000001011101001",33064 => "0000001011101000",
33065 => "0000001011100111",33066 => "0000001011100110",
33067 => "0000001011100110",33068 => "0000001011100101",
33069 => "0000000001001010",33070 => "0000001011100011",
33071 => "0000001011100011",33072 => "0000001011100010",
33073 => "0000001011100001",33074 => "0000001011100000",
33075 => "0000001011100000",33076 => "0000001011011111",
33077 => "0000001011011110",33078 => "0000001011011101",
33079 => "0000001011011101",33080 => "0000001011011100",
33081 => "0000001011011011",33082 => "0000001011011011",
33083 => "0000000001001001",33084 => "0000001011011001",
33085 => "0000001011011000",33086 => "0000001011011000",
33087 => "0000001011010111",33088 => "0000001011010110",
33089 => "0000001011010101",33090 => "0000001011010101",
33091 => "0000001011010100",33092 => "0000001011010011",
33093 => "0000001011010011",33094 => "0000001011010010",
33095 => "0000001011010001",33096 => "0000000001001000",
33097 => "0000000001001000",33098 => "0000001011001111",
33099 => "0000001011001110",33100 => "0000001011001101",
33101 => "0000001011001101",33102 => "0000001011001100",
33103 => "0000001011001011",33104 => "0000001011001011",
33105 => "0000001011001010",33106 => "0000001011001001",
33107 => "0000001011001000",33108 => "0000001011001000",
33109 => "0000001011000111",33110 => "0000000001000111",
33111 => "0000000001000111",33112 => "0000001011000101",
33113 => "0000001011000100",33114 => "0000001011000100",
33115 => "0000001011000011",33116 => "0000001011000010",
33117 => "0000001011000001",33118 => "0000001011000001",
33119 => "0000001011000000",33120 => "0000001010111111",
33121 => "0000001010111111",33122 => "0000001010111110",
33123 => "0000001010111101",33124 => "0000000000000111",
33125 => "0000000000000111",33126 => "0000001010111011",
33127 => "0000001010111010",33128 => "0000001010111010",
33129 => "0000001010111001",33130 => "0000001010111000",
33131 => "0000001010111000",33132 => "0000001010110111",
33133 => "0000001010110110",33134 => "0000001010110110",
33135 => "0000001010110101",33136 => "0000001010110100",
33137 => "0000001010110011",33138 => "0000001010110011",
33139 => "0000000001000101",33140 => "0000001010110001",
33141 => "0000001010110001",33142 => "0000001010110000",
33143 => "0000001010101111",33144 => "0000001010101111",
33145 => "0000001010101110",33146 => "0000001010101101",
33147 => "0000001010101101",33148 => "0000001010101100",
33149 => "0000001010101011",33150 => "0000001010101010",
33151 => "0000001010101010",33152 => "0000001010101001",
33153 => "0000000001000100",33154 => "0000000001000100",
33155 => "0000001010100111",33156 => "0000001010100110",
33157 => "0000001010100110",33158 => "0000001010100101",
33159 => "0000001010100100",33160 => "0000001010100100",
33161 => "0000001010100011",33162 => "0000001010100010",
33163 => "0000001010100010",33164 => "0000001010100001",
33165 => "0000001010100000",33166 => "0000001010100000",
33167 => "0000001010011111",33168 => "0000000001000011",
33169 => "0000000001000011",33170 => "0000001010011101",
33171 => "0000001010011100",33172 => "0000001010011100",
33173 => "0000001010011011",33174 => "0000001010011010",
33175 => "0000001010011010",33176 => "0000001010011001",
33177 => "0000001010011000",33178 => "0000001010011000",
33179 => "0000001010010111",33180 => "0000001010010110",
33181 => "0000001010010110",33182 => "0000001010010101",
33183 => "0000000001000010",33184 => "0000000001000010",
33185 => "0000001010010011",33186 => "0000001010010010",
33187 => "0000001010010010",33188 => "0000001010010001",
33189 => "0000001010010000",33190 => "0000001010010000",
33191 => "0000001010001111",33192 => "0000001010001110",
33193 => "0000001010001110",33194 => "0000001010001101",
33195 => "0000001010001100",33196 => "0000001010001100",
33197 => "0000001010001011",33198 => "0000001010001011",
33199 => "0000000001000001",33200 => "0000001010001001",
33201 => "0000001010001001",33202 => "0000001010001000",
33203 => "0000001010000111",33204 => "0000001010000111",
33205 => "0000001010000110",33206 => "0000001010000101",
33207 => "0000001010000101",33208 => "0000001010000100",
33209 => "0000001010000011",33210 => "0000001010000011",
33211 => "0000001010000010",33212 => "0000001010000001",
33213 => "0000001010000001",33214 => "0000000001000000",
33215 => "0000000001000000",33216 => "0000001001111111",
33217 => "0000001001111110",33218 => "0000001001111110",
33219 => "0000001001111101",33220 => "0000001001111100",
33221 => "0000001001111100",33222 => "0000001001111011",
33223 => "0000001001111010",33224 => "0000001001111010",
33225 => "0000001001111001",33226 => "0000001001111001",
33227 => "0000001001111000",33228 => "0000001001110111",
33229 => "0000001001110111",33230 => "0000000000111111",
33231 => "0000001001110101",33232 => "0000001001110101",
33233 => "0000001001110100",33234 => "0000001001110100",
33235 => "0000001001110011",33236 => "0000001001110010",
33237 => "0000001001110010",33238 => "0000001001110001",
33239 => "0000001001110000",33240 => "0000001001110000",
33241 => "0000001001101111",33242 => "0000001001101111",
33243 => "0000001001101110",33244 => "0000001001101101",
33245 => "0000001001101101",33246 => "0000000000111110",
33247 => "0000001001101011",33248 => "0000001001101011",
33249 => "0000001001101010",33250 => "0000001001101010",
33251 => "0000001001101001",33252 => "0000001001101000",
33253 => "0000001001101000",33254 => "0000001001100111",
33255 => "0000001001100110",33256 => "0000001001100110",
33257 => "0000001001100101",33258 => "0000001001100101",
33259 => "0000001001100100",33260 => "0000001001100011",
33261 => "0000001001100011",33262 => "0000000000111101",
33263 => "0000000000111101",33264 => "0000001001100001",
33265 => "0000001001100000",33266 => "0000001001100000",
33267 => "0000001001011111",33268 => "0000001001011111",
33269 => "0000001001011110",33270 => "0000001001011101",
33271 => "0000001001011101",33272 => "0000001001011100",
33273 => "0000001001011100",33274 => "0000001001011011",
33275 => "0000001001011010",33276 => "0000001001011010",
33277 => "0000001001011001",33278 => "0000000000000110",
33279 => "0000000000000110",33280 => "0000001001010111",
33281 => "0000001001010111",33282 => "0000001001010110",
33283 => "0000001001010110",33284 => "0000001001010101",
33285 => "0000001001010100",33286 => "0000001001010100",
33287 => "0000001001010011",33288 => "0000001001010011",
33289 => "0000001001010010",33290 => "0000001001010001",
33291 => "0000001001010001",33292 => "0000001001010000",
33293 => "0000001001010000",33294 => "0000001001001111",
33295 => "0000000000111011",33296 => "0000000000111011",
33297 => "0000001001001101",33298 => "0000001001001101",
33299 => "0000001001001100",33300 => "0000001001001011",
33301 => "0000001001001011",33302 => "0000001001001010",
33303 => "0000001001001010",33304 => "0000001001001001",
33305 => "0000001001001000",33306 => "0000001001001000",
33307 => "0000001001000111",33308 => "0000001001000111",
33309 => "0000001001000110",33310 => "0000001001000110",
33311 => "0000001001000101",33312 => "0000000000111010",
33313 => "0000000000111010",33314 => "0000001001000011",
33315 => "0000001001000011",33316 => "0000001001000010",
33317 => "0000001001000010",33318 => "0000001001000001",
33319 => "0000001001000000",33320 => "0000001001000000",
33321 => "0000001000111111",33322 => "0000001000111111",
33323 => "0000001000111110",33324 => "0000001000111101",
33325 => "0000001000111101",33326 => "0000001000111100",
33327 => "0000001000111100",33328 => "0000001000111011",
33329 => "0000001000111011",33330 => "0000000000111001",
33331 => "0000001000111001",33332 => "0000001000111001",
33333 => "0000001000111000",33334 => "0000001000111000",
33335 => "0000001000110111",33336 => "0000001000110111",
33337 => "0000001000110110",33338 => "0000001000110110",
33339 => "0000001000110101",33340 => "0000001000110100",
33341 => "0000001000110100",33342 => "0000001000110011",
33343 => "0000001000110011",33344 => "0000001000110010",
33345 => "0000001000110010",33346 => "0000001000110001",
33347 => "0000000000111000",33348 => "0000000000111000",
33349 => "0000001000101111",33350 => "0000001000101111",
33351 => "0000001000101110",33352 => "0000001000101110",
33353 => "0000001000101101",33354 => "0000001000101101",
33355 => "0000001000101100",33356 => "0000001000101011",
33357 => "0000001000101011",33358 => "0000001000101010",
33359 => "0000001000101010",33360 => "0000001000101001",
33361 => "0000001000101001",33362 => "0000001000101000",
33363 => "0000001000101000",33364 => "0000001000100111",
33365 => "0000000000110111",33366 => "0000000000110111",
33367 => "0000001000100101",33368 => "0000001000100101",
33369 => "0000001000100100",33370 => "0000001000100100",
33371 => "0000001000100011",33372 => "0000001000100011",
33373 => "0000001000100010",33374 => "0000001000100010",
33375 => "0000001000100001",33376 => "0000001000100000",
33377 => "0000001000100000",33378 => "0000001000011111",
33379 => "0000001000011111",33380 => "0000001000011110",
33381 => "0000001000011110",33382 => "0000001000011101",
33383 => "0000001000011101",33384 => "0000000000110110",
33385 => "0000000000110110",33386 => "0000001000011011",
33387 => "0000001000011010",33388 => "0000001000011010",
33389 => "0000001000011001",33390 => "0000001000011001",
33391 => "0000001000011000",33392 => "0000001000011000",
33393 => "0000001000010111",33394 => "0000001000010111",
33395 => "0000001000010110",33396 => "0000001000010110",
33397 => "0000001000010101",33398 => "0000001000010101",
33399 => "0000001000010100",33400 => "0000001000010100",
33401 => "0000001000010011",33402 => "0000000000110101",
33403 => "0000000000110101",33404 => "0000001000010001",
33405 => "0000001000010001",33406 => "0000001000010000",
33407 => "0000001000010000",33408 => "0000001000001111",
33409 => "0000001000001111",33410 => "0000001000001110",
33411 => "0000001000001110",33412 => "0000001000001101",
33413 => "0000001000001101",33414 => "0000001000001100",
33415 => "0000001000001100",33416 => "0000001000001011",
33417 => "0000001000001011",33418 => "0000001000001010",
33419 => "0000001000001010",33420 => "0000001000001001",
33421 => "0000000000110100",33422 => "0000000000110100",
33423 => "0000001000000111",33424 => "0000001000000111",
33425 => "0000001000000110",33426 => "0000001000000110",
33427 => "0000001000000101",33428 => "0000001000000101",
33429 => "0000001000000100",33430 => "0000001000000100",
33431 => "0000001000000011",33432 => "0000001000000011",
33433 => "0000001000000010",33434 => "0000001000000010",
33435 => "0000001000000001",33436 => "0000001000000001",
33437 => "0000001000000000",33438 => "0000001000000000",
33439 => "0000000111111111",33440 => "0000000111111111",
33441 => "0000000000110011",33442 => "0000000000110011",
33443 => "0000000111111101",33444 => "0000000111111101",
33445 => "0000000111111100",33446 => "0000000111111100",
33447 => "0000000111111011",33448 => "0000000111111011",
33449 => "0000000111111010",33450 => "0000000111111010",
33451 => "0000000111111001",33452 => "0000000111111001",
33453 => "0000000111111000",33454 => "0000000111111000",
33455 => "0000000111110111",33456 => "0000000111110111",
33457 => "0000000111110110",33458 => "0000000111110110",
33459 => "0000000111110101",33460 => "0000000111110101",
33461 => "0000000000000101",33462 => "0000000000000101",
33463 => "0000000111110011",33464 => "0000000111110011",
33465 => "0000000111110010",33466 => "0000000111110010",
33467 => "0000000111110001",33468 => "0000000111110001",
33469 => "0000000111110000",33470 => "0000000111110000",
33471 => "0000000111101111",33472 => "0000000111101111",
33473 => "0000000111101110",33474 => "0000000111101110",
33475 => "0000000111101101",33476 => "0000000111101101",
33477 => "0000000111101100",33478 => "0000000111101100",
33479 => "0000000111101011",33480 => "0000000111101011",
33481 => "0000000000110001",33482 => "0000000000110001",
33483 => "0000000111101001",33484 => "0000000111101001",
33485 => "0000000111101000",33486 => "0000000111101000",
33487 => "0000000111100111",33488 => "0000000111100111",
33489 => "0000000111100110",33490 => "0000000111100110",
33491 => "0000000111100101",33492 => "0000000111100101",
33493 => "0000000111100100",33494 => "0000000111100100",
33495 => "0000000111100011",33496 => "0000000111100011",
33497 => "0000000111100010",33498 => "0000000111100010",
33499 => "0000000111100001",33500 => "0000000111100001",
33501 => "0000000000110000",33502 => "0000000000110000",
33503 => "0000000000110000",33504 => "0000000111011111",
33505 => "0000000111011111",33506 => "0000000111011110",
33507 => "0000000111011110",33508 => "0000000111011101",
33509 => "0000000111011101",33510 => "0000000111011100",
33511 => "0000000111011100",33512 => "0000000111011011",
33513 => "0000000111011011",33514 => "0000000111011010",
33515 => "0000000111011010",33516 => "0000000111011001",
33517 => "0000000111011001",33518 => "0000000111011000",
33519 => "0000000111011000",33520 => "0000000111010111",
33521 => "0000000111010111",33522 => "0000000000101111",
33523 => "0000000000101111",33524 => "0000000000101111",
33525 => "0000000111010101",33526 => "0000000111010101",
33527 => "0000000111010100",33528 => "0000000111010100",
33529 => "0000000111010011",33530 => "0000000111010011",
33531 => "0000000111010010",33532 => "0000000111010010",
33533 => "0000000111010001",33534 => "0000000111010001",
33535 => "0000000111010000",33536 => "0000000111010000",
33537 => "0000000111001111",33538 => "0000000111001111",
33539 => "0000000111001111",33540 => "0000000111001110",
33541 => "0000000111001110",33542 => "0000000111001101",
33543 => "0000000111001101",33544 => "0000000000101110",
33545 => "0000000000101110",33546 => "0000000111001011",
33547 => "0000000111001011",33548 => "0000000111001010",
33549 => "0000000111001010",33550 => "0000000111001001",
33551 => "0000000111001001",33552 => "0000000111001001",
33553 => "0000000111001000",33554 => "0000000111001000",
33555 => "0000000111000111",33556 => "0000000111000111",
33557 => "0000000111000110",33558 => "0000000111000110",
33559 => "0000000111000101",33560 => "0000000111000101",
33561 => "0000000111000100",33562 => "0000000111000100",
33563 => "0000000111000100",33564 => "0000000111000011",
33565 => "0000000111000011",33566 => "0000000000101101",
33567 => "0000000000101101",33568 => "0000000111000001",
33569 => "0000000111000001",33570 => "0000000111000000",
33571 => "0000000111000000",33572 => "0000000111000000",
33573 => "0000000110111111",33574 => "0000000110111111",
33575 => "0000000110111110",33576 => "0000000110111110",
33577 => "0000000110111101",33578 => "0000000110111101",
33579 => "0000000110111100",33580 => "0000000110111100",
33581 => "0000000110111100",33582 => "0000000110111011",
33583 => "0000000110111011",33584 => "0000000110111010",
33585 => "0000000110111010",33586 => "0000000110111001",
33587 => "0000000110111001",33588 => "0000000000101100",
33589 => "0000000000101100",33590 => "0000000000101100",
33591 => "0000000110110111",33592 => "0000000110110111",
33593 => "0000000110110110",33594 => "0000000110110110",
33595 => "0000000110110101",33596 => "0000000110110101",
33597 => "0000000110110100",33598 => "0000000110110100",
33599 => "0000000110110100",33600 => "0000000110110011",
33601 => "0000000110110011",33602 => "0000000110110010",
33603 => "0000000110110010",33604 => "0000000110110001",
33605 => "0000000110110001",33606 => "0000000110110001",
33607 => "0000000110110000",33608 => "0000000110110000",
33609 => "0000000110101111",33610 => "0000000110101111",
33611 => "0000000000101011",33612 => "0000000000101011",
33613 => "0000000000101011",33614 => "0000000110101101",
33615 => "0000000110101101",33616 => "0000000110101100",
33617 => "0000000110101100",33618 => "0000000110101011",
33619 => "0000000110101011",33620 => "0000000110101011",
33621 => "0000000110101010",33622 => "0000000110101010",
33623 => "0000000110101001",33624 => "0000000110101001",
33625 => "0000000110101000",33626 => "0000000110101000",
33627 => "0000000110101000",33628 => "0000000110100111",
33629 => "0000000110100111",33630 => "0000000110100110",
33631 => "0000000110100110",33632 => "0000000110100101",
33633 => "0000000110100101",33634 => "0000000110100101",
33635 => "0000000000101010",33636 => "0000000000101010",
33637 => "0000000110100011",33638 => "0000000110100011",
33639 => "0000000110100011",33640 => "0000000110100010",
33641 => "0000000110100010",33642 => "0000000110100001",
33643 => "0000000110100001",33644 => "0000000110100000",
33645 => "0000000110100000",33646 => "0000000110100000",
33647 => "0000000110011111",33648 => "0000000110011111",
33649 => "0000000110011110",33650 => "0000000110011110",
33651 => "0000000110011110",33652 => "0000000110011101",
33653 => "0000000110011101",33654 => "0000000110011100",
33655 => "0000000110011100",33656 => "0000000110011011",
33657 => "0000000110011011",33658 => "0000000110011011",
33659 => "0000000000101001",33660 => "0000000000101001",
33661 => "0000000110011001",33662 => "0000000110011001",
33663 => "0000000110011001",33664 => "0000000110011000",
33665 => "0000000110011000",33666 => "0000000110010111",
33667 => "0000000110010111",33668 => "0000000110010111",
33669 => "0000000110010110",33670 => "0000000110010110",
33671 => "0000000110010101",33672 => "0000000110010101",
33673 => "0000000110010101",33674 => "0000000110010100",
33675 => "0000000110010100",33676 => "0000000110010011",
33677 => "0000000110010011",33678 => "0000000110010011",
33679 => "0000000110010010",33680 => "0000000110010010",
33681 => "0000000110010001",33682 => "0000000110010001",
33683 => "0000000110010001",33684 => "0000000000000100",
33685 => "0000000000000100",33686 => "0000000110001111",
33687 => "0000000110001111",33688 => "0000000110001111",
33689 => "0000000110001110",33690 => "0000000110001110",
33691 => "0000000110001101",33692 => "0000000110001101",
33693 => "0000000110001101",33694 => "0000000110001100",
33695 => "0000000110001100",33696 => "0000000110001011",
33697 => "0000000110001011",33698 => "0000000110001011",
33699 => "0000000110001010",33700 => "0000000110001010",
33701 => "0000000110001001",33702 => "0000000110001001",
33703 => "0000000110001001",33704 => "0000000110001000",
33705 => "0000000110001000",33706 => "0000000110000111",
33707 => "0000000110000111",33708 => "0000000110000111",
33709 => "0000000000100111",33710 => "0000000000100111",
33711 => "0000000110000101",33712 => "0000000110000101",
33713 => "0000000110000101",33714 => "0000000110000100",
33715 => "0000000110000100",33716 => "0000000110000100",
33717 => "0000000110000011",33718 => "0000000110000011",
33719 => "0000000110000010",33720 => "0000000110000010",
33721 => "0000000110000010",33722 => "0000000110000001",
33723 => "0000000110000001",33724 => "0000000110000000",
33725 => "0000000110000000",33726 => "0000000110000000",
33727 => "0000000101111111",33728 => "0000000101111111",
33729 => "0000000101111111",33730 => "0000000101111110",
33731 => "0000000101111110",33732 => "0000000101111101",
33733 => "0000000101111101",33734 => "0000000101111101",
33735 => "0000000000100110",33736 => "0000000000100110",
33737 => "0000000101111011",33738 => "0000000101111011",
33739 => "0000000101111011",33740 => "0000000101111010",
33741 => "0000000101111010",33742 => "0000000101111010",
33743 => "0000000101111001",33744 => "0000000101111001",
33745 => "0000000101111000",33746 => "0000000101111000",
33747 => "0000000101111000",33748 => "0000000101110111",
33749 => "0000000101110111",33750 => "0000000101110111",
33751 => "0000000101110110",33752 => "0000000101110110",
33753 => "0000000101110101",33754 => "0000000101110101",
33755 => "0000000101110101",33756 => "0000000101110100",
33757 => "0000000101110100",33758 => "0000000101110100",
33759 => "0000000101110011",33760 => "0000000101110011",
33761 => "0000000000100101",33762 => "0000000000100101",
33763 => "0000000000100101",33764 => "0000000101110001",
33765 => "0000000101110001",33766 => "0000000101110001",
33767 => "0000000101110000",33768 => "0000001110001001",
33769 => "0000001110001001",33770 => "0000001110001001",
33771 => "0000001110001001",33772 => "0000001110001000",
33773 => "0000001110001000",33774 => "0000001110001000",
33775 => "0000001110001000",33776 => "0000001110001000",
33777 => "0000001110001000",33778 => "0000001110001000",
33779 => "0000001110001000",33780 => "0000001110001000",
33781 => "0000001110001000",33782 => "0000001110001000",
33783 => "0000001110000111",33784 => "0000001110000111",
33785 => "0000001110000111",33786 => "0000001110000111",
33787 => "0000001110000111",33788 => "0000001110000111",
33789 => "0000001110000111",33790 => "0000001110000111",
33791 => "0000001110000111",33792 => "0000001110000111",
33793 => "0000001110000111",33794 => "0000001110000110",
33795 => "0000001110000110",33796 => "0000001110000110",
33797 => "0000001110000110",33798 => "0000001110000110",
33799 => "0000001110000110",33800 => "0000001110000110",
33801 => "0000001110000110",33802 => "0000001110000110",
33803 => "0000001110000110",33804 => "0000001110000110",
33805 => "0000001110000101",33806 => "0000001110000101",
33807 => "0000001110000101",33808 => "0000001110000101",
33809 => "0000001110000101",33810 => "0000001110000101",
33811 => "0000001110000101",33812 => "0000001110000101",
33813 => "0000001110000101",33814 => "0000001110000101",
33815 => "0000001110000101",33816 => "0000001110000101",
33817 => "0000000000001001",33818 => "0000000000001001",
33819 => "0000000000001001",33820 => "0000000000001001",
33821 => "0000000000001001",33822 => "0000000000001001",
33823 => "0000000000001001",33824 => "0000000000001001",
33825 => "0000000000001001",33826 => "0000000000001001",
33827 => "0000000000001001",33828 => "0000001110000011",
33829 => "0000001110000011",33830 => "0000001110000011",
33831 => "0000001110000011",33832 => "0000001110000011",
33833 => "0000001110000011",33834 => "0000001110000011",
33835 => "0000001110000011",33836 => "0000001110000011",
33837 => "0000001110000011",33838 => "0000001110000011",
33839 => "0000001110000010",33840 => "0000001110000010",
33841 => "0000001110000010",33842 => "0000001110000010",
33843 => "0000001110000010",33844 => "0000001110000010",
33845 => "0000001110000010",33846 => "0000001110000010",
33847 => "0000001110000010",33848 => "0000001110000010",
33849 => "0000001110000010",33850 => "0000001110000001",
33851 => "0000001110000001",33852 => "0000001110000001",
33853 => "0000001110000001",33854 => "0000001110000001",
33855 => "0000001110000001",33856 => "0000001110000001",
33857 => "0000001110000001",33858 => "0000001110000001",
33859 => "0000001110000001",33860 => "0000001110000001",
33861 => "0000001110000000",33862 => "0000001110000000",
33863 => "0000001110000000",33864 => "0000001110000000",
33865 => "0000001110000000",33866 => "0000001110000000",
33867 => "0000001110000000",33868 => "0000001110000000",
33869 => "0000001110000000",33870 => "0000001110000000",
33871 => "0000001110000000",33872 => "0000001101111111",
33873 => "0000001101111111",33874 => "0000001101111111",
33875 => "0000001101111111",33876 => "0000001101111111",
33877 => "0000001101111111",33878 => "0000001101111111",
33879 => "0000001101111111",33880 => "0000001101111111",
33881 => "0000001101111111",33882 => "0000001101111111",
33883 => "0000001101111110",33884 => "0000001101111110",
33885 => "0000001101111110",33886 => "0000001101111110",
33887 => "0000001101111110",33888 => "0000001101111110",
33889 => "0000001101111110",33890 => "0000001101111110",
33891 => "0000001101111110",33892 => "0000001101111110",
33893 => "0000001101111110",33894 => "0000001101111110",
33895 => "0000001101111101",33896 => "0000001101111101",
33897 => "0000001101111101",33898 => "0000001101111101",
33899 => "0000001101111101",33900 => "0000001101111101",
33901 => "0000001101111101",33902 => "0000001101111101",
33903 => "0000001101111101",33904 => "0000001101111101",
33905 => "0000001101111101",33906 => "0000001101111100",
33907 => "0000001101111100",33908 => "0000001101111100",
33909 => "0000001101111100",33910 => "0000001101111100",
33911 => "0000001101111100",33912 => "0000001101111100",
33913 => "0000001101111100",33914 => "0000001101111100",
33915 => "0000001101111100",33916 => "0000001101111100",
33917 => "0000001101111011",33918 => "0000001101111011",
33919 => "0000001101111011",33920 => "0000001101111011",
33921 => "0000001101111011",33922 => "0000001101111011",
33923 => "0000001101111011",33924 => "0000001101111011",
33925 => "0000001101111011",33926 => "0000001101111011",
33927 => "0000001101111011",33928 => "0000000001011001",
33929 => "0000000001011001",33930 => "0000000001011001",
33931 => "0000000001011001",33932 => "0000000001011001",
33933 => "0000000001011001",33934 => "0000000001011001",
33935 => "0000000001011001",33936 => "0000000001011001",
33937 => "0000000001011001",33938 => "0000000001011001",
33939 => "0000001101111001",33940 => "0000001101111001",
33941 => "0000001101111001",33942 => "0000001101111001",
33943 => "0000001101111001",33944 => "0000001101111001",
33945 => "0000001101111001",33946 => "0000001101111001",
33947 => "0000001101111001",33948 => "0000001101111001",
33949 => "0000001101111001",33950 => "0000001101111001",
33951 => "0000001101111000",33952 => "0000001101111000",
33953 => "0000001101111000",33954 => "0000001101111000",
33955 => "0000001101111000",33956 => "0000001101111000",
33957 => "0000001101111000",33958 => "0000001101111000",
33959 => "0000001101111000",33960 => "0000001101111000",
33961 => "0000001101111000",33962 => "0000001101110111",
33963 => "0000001101110111",33964 => "0000001101110111",
33965 => "0000001101110111",33966 => "0000001101110111",
33967 => "0000001101110111",33968 => "0000001101110111",
33969 => "0000001101110111",33970 => "0000001101110111",
33971 => "0000001101110111",33972 => "0000001101110111",
33973 => "0000001101110110",33974 => "0000001101110110",
33975 => "0000001101110110",33976 => "0000001101110110",
33977 => "0000001101110110",33978 => "0000001101110110",
33979 => "0000001101110110",33980 => "0000001101110110",
33981 => "0000001101110110",33982 => "0000001101110110",
33983 => "0000001101110110",33984 => "0000001101110110",
33985 => "0000001101110101",33986 => "0000001101110101",
33987 => "0000001101110101",33988 => "0000001101110101",
33989 => "0000001101110101",33990 => "0000001101110101",
33991 => "0000001101110101",33992 => "0000001101110101",
33993 => "0000001101110101",33994 => "0000001101110101",
33995 => "0000001101110101",33996 => "0000001101110100",
33997 => "0000001101110100",33998 => "0000001101110100",
33999 => "0000001101110100",34000 => "0000001101110100",
34001 => "0000001101110100",34002 => "0000001101110100",
34003 => "0000001101110100",34004 => "0000001101110100",
34005 => "0000001101110100",34006 => "0000001101110100",
34007 => "0000001101110011",34008 => "0000001101110011",
34009 => "0000001101110011",34010 => "0000001101110011",
34011 => "0000001101110011",34012 => "0000001101110011",
34013 => "0000001101110011",34014 => "0000001101110011",
34015 => "0000001101110011",34016 => "0000001101110011",
34017 => "0000001101110011",34018 => "0000001101110010",
34019 => "0000001101110010",34020 => "0000001101110010",
34021 => "0000001101110010",34022 => "0000001101110010",
34023 => "0000001101110010",34024 => "0000001101110010",
34025 => "0000001101110010",34026 => "0000001101110010",
34027 => "0000001101110010",34028 => "0000001101110010",
34029 => "0000001101110010",34030 => "0000001101110001",
34031 => "0000001101110001",34032 => "0000001101110001",
34033 => "0000001101110001",34034 => "0000001101110001",
34035 => "0000001101110001",34036 => "0000001101110001",
34037 => "0000001101110001",34038 => "0000001101110001",
34039 => "0000001101110001",34040 => "0000001101110001",
34041 => "0000000001011000",34042 => "0000000001011000",
34043 => "0000000001011000",34044 => "0000000001011000",
34045 => "0000000001011000",34046 => "0000000001011000",
34047 => "0000000001011000",34048 => "0000000001011000",
34049 => "0000000001011000",34050 => "0000000001011000",
34051 => "0000000001011000",34052 => "0000000001011000",
34053 => "0000001101101111",34054 => "0000001101101111",
34055 => "0000001101101111",34056 => "0000001101101111",
34057 => "0000001101101111",34058 => "0000001101101111",
34059 => "0000001101101111",34060 => "0000001101101111",
34061 => "0000001101101111",34062 => "0000001101101111",
34063 => "0000001101101111",34064 => "0000001101101110",
34065 => "0000001101101110",34066 => "0000001101101110",
34067 => "0000001101101110",34068 => "0000001101101110",
34069 => "0000001101101110",34070 => "0000001101101110",
34071 => "0000001101101110",34072 => "0000001101101110",
34073 => "0000001101101110",34074 => "0000001101101110",
34075 => "0000001101101101",34076 => "0000001101101101",
34077 => "0000001101101101",34078 => "0000001101101101",
34079 => "0000001101101101",34080 => "0000001101101101",
34081 => "0000001101101101",34082 => "0000001101101101",
34083 => "0000001101101101",34084 => "0000001101101101",
34085 => "0000001101101101",34086 => "0000001101101101",
34087 => "0000001101101100",34088 => "0000001101101100",
34089 => "0000001101101100",34090 => "0000001101101100",
34091 => "0000001101101100",34092 => "0000001101101100",
34093 => "0000001101101100",34094 => "0000001101101100",
34095 => "0000001101101100",34096 => "0000001101101100",
34097 => "0000001101101100",34098 => "0000001101101011",
34099 => "0000001101101011",34100 => "0000001101101011",
34101 => "0000001101101011",34102 => "0000001101101011",
34103 => "0000001101101011",34104 => "0000001101101011",
34105 => "0000001101101011",34106 => "0000001101101011",
34107 => "0000001101101011",34108 => "0000001101101011",
34109 => "0000001101101011",34110 => "0000001101101010",
34111 => "0000001101101010",34112 => "0000001101101010",
34113 => "0000001101101010",34114 => "0000001101101010",
34115 => "0000001101101010",34116 => "0000001101101010",
34117 => "0000001101101010",34118 => "0000001101101010",
34119 => "0000001101101010",34120 => "0000001101101010",
34121 => "0000001101101001",34122 => "0000001101101001",
34123 => "0000001101101001",34124 => "0000001101101001",
34125 => "0000001101101001",34126 => "0000001101101001",
34127 => "0000001101101001",34128 => "0000001101101001",
34129 => "0000001101101001",34130 => "0000001101101001",
34131 => "0000001101101001",34132 => "0000001101101000",
34133 => "0000001101101000",34134 => "0000001101101000",
34135 => "0000001101101000",34136 => "0000001101101000",
34137 => "0000001101101000",34138 => "0000001101101000",
34139 => "0000001101101000",34140 => "0000001101101000",
34141 => "0000001101101000",34142 => "0000001101101000",
34143 => "0000001101101000",34144 => "0000001101100111",
34145 => "0000001101100111",34146 => "0000001101100111",
34147 => "0000001101100111",34148 => "0000001101100111",
34149 => "0000001101100111",34150 => "0000001101100111",
34151 => "0000001101100111",34152 => "0000001101100111",
34153 => "0000001101100111",34154 => "0000001101100111",
34155 => "0000000001010111",34156 => "0000000001010111",
34157 => "0000000001010111",34158 => "0000000001010111",
34159 => "0000000001010111",34160 => "0000000001010111",
34161 => "0000000001010111",34162 => "0000000001010111",
34163 => "0000000001010111",34164 => "0000000001010111",
34165 => "0000000001010111",34166 => "0000000001010111",
34167 => "0000001101100101",34168 => "0000001101100101",
34169 => "0000001101100101",34170 => "0000001101100101",
34171 => "0000001101100101",34172 => "0000001101100101",
34173 => "0000001101100101",34174 => "0000001101100101",
34175 => "0000001101100101",34176 => "0000001101100101",
34177 => "0000001101100101",34178 => "0000001101100100",
34179 => "0000001101100100",34180 => "0000001101100100",
34181 => "0000001101100100",34182 => "0000001101100100",
34183 => "0000001101100100",34184 => "0000001101100100",
34185 => "0000001101100100",34186 => "0000001101100100",
34187 => "0000001101100100",34188 => "0000001101100100",
34189 => "0000001101100100",34190 => "0000001101100011",
34191 => "0000001101100011",34192 => "0000001101100011",
34193 => "0000001101100011",34194 => "0000001101100011",
34195 => "0000001101100011",34196 => "0000001101100011",
34197 => "0000001101100011",34198 => "0000001101100011",
34199 => "0000001101100011",34200 => "0000001101100011",
34201 => "0000001101100010",34202 => "0000001101100010",
34203 => "0000001101100010",34204 => "0000001101100010",
34205 => "0000001101100010",34206 => "0000001101100010",
34207 => "0000001101100010",34208 => "0000001101100010",
34209 => "0000001101100010",34210 => "0000001101100010",
34211 => "0000001101100010",34212 => "0000001101100010",
34213 => "0000001101100001",34214 => "0000001101100001",
34215 => "0000001101100001",34216 => "0000001101100001",
34217 => "0000001101100001",34218 => "0000001101100001",
34219 => "0000001101100001",34220 => "0000001101100001",
34221 => "0000001101100001",34222 => "0000001101100001",
34223 => "0000001101100001",34224 => "0000001101100001",
34225 => "0000001101100000",34226 => "0000001101100000",
34227 => "0000001101100000",34228 => "0000001101100000",
34229 => "0000001101100000",34230 => "0000001101100000",
34231 => "0000001101100000",34232 => "0000001101100000",
34233 => "0000001101100000",34234 => "0000001101100000",
34235 => "0000001101100000",34236 => "0000001101011111",
34237 => "0000001101011111",34238 => "0000001101011111",
34239 => "0000001101011111",34240 => "0000001101011111",
34241 => "0000001101011111",34242 => "0000001101011111",
34243 => "0000001101011111",34244 => "0000001101011111",
34245 => "0000001101011111",34246 => "0000001101011111",
34247 => "0000001101011111",34248 => "0000001101011110",
34249 => "0000001101011110",34250 => "0000001101011110",
34251 => "0000001101011110",34252 => "0000001101011110",
34253 => "0000001101011110",34254 => "0000001101011110",
34255 => "0000001101011110",34256 => "0000001101011110",
34257 => "0000001101011110",34258 => "0000001101011110",
34259 => "0000001101011101",34260 => "0000001101011101",
34261 => "0000001101011101",34262 => "0000001101011101",
34263 => "0000001101011101",34264 => "0000001101011101",
34265 => "0000001101011101",34266 => "0000001101011101",
34267 => "0000001101011101",34268 => "0000001101011101",
34269 => "0000001101011101",34270 => "0000001101011101",
34271 => "0000000001010110",34272 => "0000000001010110",
34273 => "0000000001010110",34274 => "0000000001010110",
34275 => "0000000001010110",34276 => "0000000001010110",
34277 => "0000000001010110",34278 => "0000000001010110",
34279 => "0000000001010110",34280 => "0000000001010110",
34281 => "0000000001010110",34282 => "0000000001010110",
34283 => "0000001101011011",34284 => "0000001101011011",
34285 => "0000001101011011",34286 => "0000001101011011",
34287 => "0000001101011011",34288 => "0000001101011011",
34289 => "0000001101011011",34290 => "0000001101011011",
34291 => "0000001101011011",34292 => "0000001101011011",
34293 => "0000001101011011",34294 => "0000001101011010",
34295 => "0000001101011010",34296 => "0000001101011010",
34297 => "0000001101011010",34298 => "0000001101011010",
34299 => "0000001101011010",34300 => "0000001101011010",
34301 => "0000001101011010",34302 => "0000001101011010",
34303 => "0000001101011010",34304 => "0000001101011010",
34305 => "0000001101011010",34306 => "0000001101011001",
34307 => "0000001101011001",34308 => "0000001101011001",
34309 => "0000001101011001",34310 => "0000001101011001",
34311 => "0000001101011001",34312 => "0000001101011001",
34313 => "0000001101011001",34314 => "0000001101011001",
34315 => "0000001101011001",34316 => "0000001101011001",
34317 => "0000001101011001",34318 => "0000001101011000",
34319 => "0000001101011000",34320 => "0000001101011000",
34321 => "0000001101011000",34322 => "0000001101011000",
34323 => "0000001101011000",34324 => "0000001101011000",
34325 => "0000001101011000",34326 => "0000001101011000",
34327 => "0000001101011000",34328 => "0000001101011000",
34329 => "0000001101010111",34330 => "0000001101010111",
34331 => "0000001101010111",34332 => "0000001101010111",
34333 => "0000001101010111",34334 => "0000001101010111",
34335 => "0000001101010111",34336 => "0000001101010111",
34337 => "0000001101010111",34338 => "0000001101010111",
34339 => "0000001101010111",34340 => "0000001101010111",
34341 => "0000001101010110",34342 => "0000001101010110",
34343 => "0000001101010110",34344 => "0000001101010110",
34345 => "0000001101010110",34346 => "0000001101010110",
34347 => "0000001101010110",34348 => "0000001101010110",
34349 => "0000001101010110",34350 => "0000001101010110",
34351 => "0000001101010110",34352 => "0000001101010110",
34353 => "0000001101010101",34354 => "0000001101010101",
34355 => "0000001101010101",34356 => "0000001101010101",
34357 => "0000001101010101",34358 => "0000001101010101",
34359 => "0000001101010101",34360 => "0000001101010101",
34361 => "0000001101010101",34362 => "0000001101010101",
34363 => "0000001101010101",34364 => "0000001101010100",
34365 => "0000001101010100",34366 => "0000001101010100",
34367 => "0000001101010100",34368 => "0000001101010100",
34369 => "0000001101010100",34370 => "0000001101010100",
34371 => "0000001101010100",34372 => "0000001101010100",
34373 => "0000001101010100",34374 => "0000001101010100",
34375 => "0000001101010100",34376 => "0000001101010011",
34377 => "0000001101010011",34378 => "0000001101010011",
34379 => "0000001101010011",34380 => "0000001101010011",
34381 => "0000001101010011",34382 => "0000001101010011",
34383 => "0000001101010011",34384 => "0000001101010011",
34385 => "0000001101010011",34386 => "0000001101010011",
34387 => "0000001101010011",34388 => "0000000001010101",
34389 => "0000000001010101",34390 => "0000000001010101",
34391 => "0000000001010101",34392 => "0000000001010101",
34393 => "0000000001010101",34394 => "0000000001010101",
34395 => "0000000001010101",34396 => "0000000001010101",
34397 => "0000000001010101",34398 => "0000000001010101",
34399 => "0000000001010101",34400 => "0000001101010001",
34401 => "0000001101010001",34402 => "0000001101010001",
34403 => "0000001101010001",34404 => "0000001101010001",
34405 => "0000001101010001",34406 => "0000001101010001",
34407 => "0000001101010001",34408 => "0000001101010001",
34409 => "0000001101010001",34410 => "0000001101010001",
34411 => "0000001101010000",34412 => "0000001101010000",
34413 => "0000001101010000",34414 => "0000001101010000",
34415 => "0000001101010000",34416 => "0000001101010000",
34417 => "0000001101010000",34418 => "0000001101010000",
34419 => "0000001101010000",34420 => "0000001101010000",
34421 => "0000001101010000",34422 => "0000001101010000",
34423 => "0000001101001111",34424 => "0000001101001111",
34425 => "0000001101001111",34426 => "0000001101001111",
34427 => "0000001101001111",34428 => "0000001101001111",
34429 => "0000001101001111",34430 => "0000001101001111",
34431 => "0000001101001111",34432 => "0000001101001111",
34433 => "0000001101001111",34434 => "0000001101001111",
34435 => "0000001101001110",34436 => "0000001101001110",
34437 => "0000001101001110",34438 => "0000001101001110",
34439 => "0000001101001110",34440 => "0000001101001110",
34441 => "0000001101001110",34442 => "0000001101001110",
34443 => "0000001101001110",34444 => "0000001101001110",
34445 => "0000001101001110",34446 => "0000001101001110",
34447 => "0000001101001101",34448 => "0000001101001101",
34449 => "0000001101001101",34450 => "0000001101001101",
34451 => "0000001101001101",34452 => "0000001101001101",
34453 => "0000001101001101",34454 => "0000001101001101",
34455 => "0000001101001101",34456 => "0000001101001101",
34457 => "0000001101001101",34458 => "0000001101001101",
34459 => "0000001101001100",34460 => "0000001101001100",
34461 => "0000001101001100",34462 => "0000001101001100",
34463 => "0000001101001100",34464 => "0000001101001100",
34465 => "0000001101001100",34466 => "0000001101001100",
34467 => "0000001101001100",34468 => "0000001101001100",
34469 => "0000001101001100",34470 => "0000001101001011",
34471 => "0000001101001011",34472 => "0000001101001011",
34473 => "0000001101001011",34474 => "0000001101001011",
34475 => "0000001101001011",34476 => "0000001101001011",
34477 => "0000001101001011",34478 => "0000001101001011",
34479 => "0000001101001011",34480 => "0000001101001011",
34481 => "0000001101001011",34482 => "0000001101001010",
34483 => "0000001101001010",34484 => "0000001101001010",
34485 => "0000001101001010",34486 => "0000001101001010",
34487 => "0000001101001010",34488 => "0000001101001010",
34489 => "0000001101001010",34490 => "0000001101001010",
34491 => "0000001101001010",34492 => "0000001101001010",
34493 => "0000001101001010",34494 => "0000001101001001",
34495 => "0000001101001001",34496 => "0000001101001001",
34497 => "0000001101001001",34498 => "0000001101001001",
34499 => "0000001101001001",34500 => "0000001101001001",
34501 => "0000001101001001",34502 => "0000001101001001",
34503 => "0000001101001001",34504 => "0000001101001001",
34505 => "0000001101001001",34506 => "0000000001010100",
34507 => "0000000001010100",34508 => "0000000001010100",
34509 => "0000000001010100",34510 => "0000000001010100",
34511 => "0000000001010100",34512 => "0000000001010100",
34513 => "0000000001010100",34514 => "0000000001010100",
34515 => "0000000001010100",34516 => "0000000001010100",
34517 => "0000000001010100",34518 => "0000001101000111",
34519 => "0000001101000111",34520 => "0000001101000111",
34521 => "0000001101000111",34522 => "0000001101000111",
34523 => "0000001101000111",34524 => "0000001101000111",
34525 => "0000001101000111",34526 => "0000001101000111",
34527 => "0000001101000111",34528 => "0000001101000111",
34529 => "0000001101000111",34530 => "0000001101000110",
34531 => "0000001101000110",34532 => "0000001101000110",
34533 => "0000001101000110",34534 => "0000001101000110",
34535 => "0000001101000110",34536 => "0000001101000110",
34537 => "0000001101000110",34538 => "0000001101000110",
34539 => "0000001101000110",34540 => "0000001101000110",
34541 => "0000001101000110",34542 => "0000001101000101",
34543 => "0000001101000101",34544 => "0000001101000101",
34545 => "0000001101000101",34546 => "0000001101000101",
34547 => "0000001101000101",34548 => "0000001101000101",
34549 => "0000001101000101",34550 => "0000001101000101",
34551 => "0000001101000101",34552 => "0000001101000101",
34553 => "0000001101000101",34554 => "0000001101000100",
34555 => "0000001101000100",34556 => "0000001101000100",
34557 => "0000001101000100",34558 => "0000001101000100",
34559 => "0000001101000100",34560 => "0000001101000100",
34561 => "0000001101000100",34562 => "0000001101000100",
34563 => "0000001101000100",34564 => "0000001101000100",
34565 => "0000001101000100",34566 => "0000001101000011",
34567 => "0000001101000011",34568 => "0000001101000011",
34569 => "0000001101000011",34570 => "0000001101000011",
34571 => "0000001101000011",34572 => "0000001101000011",
34573 => "0000001101000011",34574 => "0000001101000011",
34575 => "0000001101000011",34576 => "0000001101000011",
34577 => "0000001101000011",34578 => "0000001101000010",
34579 => "0000001101000010",34580 => "0000001101000010",
34581 => "0000001101000010",34582 => "0000001101000010",
34583 => "0000001101000010",34584 => "0000001101000010",
34585 => "0000001101000010",34586 => "0000001101000010",
34587 => "0000001101000010",34588 => "0000001101000010",
34589 => "0000001101000010",34590 => "0000001101000001",
34591 => "0000001101000001",34592 => "0000001101000001",
34593 => "0000001101000001",34594 => "0000001101000001",
34595 => "0000001101000001",34596 => "0000001101000001",
34597 => "0000001101000001",34598 => "0000001101000001",
34599 => "0000001101000001",34600 => "0000001101000001",
34601 => "0000001101000001",34602 => "0000001101000000",
34603 => "0000001101000000",34604 => "0000001101000000",
34605 => "0000001101000000",34606 => "0000001101000000",
34607 => "0000001101000000",34608 => "0000001101000000",
34609 => "0000001101000000",34610 => "0000001101000000",
34611 => "0000001101000000",34612 => "0000001101000000",
34613 => "0000001101000000",34614 => "0000001100111111",
34615 => "0000001100111111",34616 => "0000001100111111",
34617 => "0000001100111111",34618 => "0000001100111111",
34619 => "0000001100111111",34620 => "0000001100111111",
34621 => "0000001100111111",34622 => "0000001100111111",
34623 => "0000001100111111",34624 => "0000001100111111",
34625 => "0000001100111111",34626 => "0000000001010011",
34627 => "0000000001010011",34628 => "0000000001010011",
34629 => "0000000001010011",34630 => "0000000001010011",
34631 => "0000000001010011",34632 => "0000000001010011",
34633 => "0000000001010011",34634 => "0000000001010011",
34635 => "0000000001010011",34636 => "0000000001010011",
34637 => "0000000001010011",34638 => "0000001100111101",
34639 => "0000001100111101",34640 => "0000001100111101",
34641 => "0000001100111101",34642 => "0000001100111101",
34643 => "0000001100111101",34644 => "0000001100111101",
34645 => "0000001100111101",34646 => "0000001100111101",
34647 => "0000001100111101",34648 => "0000001100111101",
34649 => "0000001100111101",34650 => "0000001100111100",
34651 => "0000001100111100",34652 => "0000001100111100",
34653 => "0000001100111100",34654 => "0000001100111100",
34655 => "0000001100111100",34656 => "0000001100111100",
34657 => "0000001100111100",34658 => "0000001100111100",
34659 => "0000001100111100",34660 => "0000001100111100",
34661 => "0000001100111100",34662 => "0000001100111011",
34663 => "0000001100111011",34664 => "0000001100111011",
34665 => "0000001100111011",34666 => "0000001100111011",
34667 => "0000001100111011",34668 => "0000001100111011",
34669 => "0000001100111011",34670 => "0000001100111011",
34671 => "0000001100111011",34672 => "0000001100111011",
34673 => "0000001100111011",34674 => "0000001100111010",
34675 => "0000001100111010",34676 => "0000001100111010",
34677 => "0000001100111010",34678 => "0000001100111010",
34679 => "0000001100111010",34680 => "0000001100111010",
34681 => "0000001100111010",34682 => "0000001100111010",
34683 => "0000001100111010",34684 => "0000001100111010",
34685 => "0000001100111010",34686 => "0000001100111001",
34687 => "0000001100111001",34688 => "0000001100111001",
34689 => "0000001100111001",34690 => "0000001100111001",
34691 => "0000001100111001",34692 => "0000001100111001",
34693 => "0000001100111001",34694 => "0000001100111001",
34695 => "0000001100111001",34696 => "0000001100111001",
34697 => "0000001100111001",34698 => "0000001100111000",
34699 => "0000001100111000",34700 => "0000001100111000",
34701 => "0000001100111000",34702 => "0000001100111000",
34703 => "0000001100111000",34704 => "0000001100111000",
34705 => "0000001100111000",34706 => "0000001100111000",
34707 => "0000001100111000",34708 => "0000001100111000",
34709 => "0000001100111000",34710 => "0000001100110111",
34711 => "0000001100110111",34712 => "0000001100110111",
34713 => "0000001100110111",34714 => "0000001100110111",
34715 => "0000001100110111",34716 => "0000001100110111",
34717 => "0000001100110111",34718 => "0000001100110111",
34719 => "0000001100110111",34720 => "0000001100110111",
34721 => "0000001100110111",34722 => "0000001100110111",
34723 => "0000001100110110",34724 => "0000001100110110",
34725 => "0000001100110110",34726 => "0000001100110110",
34727 => "0000001100110110",34728 => "0000001100110110",
34729 => "0000001100110110",34730 => "0000001100110110",
34731 => "0000001100110110",34732 => "0000001100110110",
34733 => "0000001100110110",34734 => "0000001100110110",
34735 => "0000001100110101",34736 => "0000001100110101",
34737 => "0000001100110101",34738 => "0000001100110101",
34739 => "0000001100110101",34740 => "0000001100110101",
34741 => "0000001100110101",34742 => "0000001100110101",
34743 => "0000001100110101",34744 => "0000001100110101",
34745 => "0000001100110101",34746 => "0000001100110101",
34747 => "0000000001010010",34748 => "0000000001010010",
34749 => "0000000001010010",34750 => "0000000001010010",
34751 => "0000000001010010",34752 => "0000000001010010",
34753 => "0000000001010010",34754 => "0000000001010010",
34755 => "0000000001010010",34756 => "0000000001010010",
34757 => "0000000001010010",34758 => "0000000001010010",
34759 => "0000001100110011",34760 => "0000001100110011",
34761 => "0000001100110011",34762 => "0000001100110011",
34763 => "0000001100110011",34764 => "0000001100110011",
34765 => "0000001100110011",34766 => "0000001100110011",
34767 => "0000001100110011",34768 => "0000001100110011",
34769 => "0000001100110011",34770 => "0000001100110011",
34771 => "0000001100110010",34772 => "0000001100110010",
34773 => "0000001100110010",34774 => "0000001100110010",
34775 => "0000001100110010",34776 => "0000001100110010",
34777 => "0000001100110010",34778 => "0000001100110010",
34779 => "0000001100110010",34780 => "0000001100110010",
34781 => "0000001100110010",34782 => "0000001100110010",
34783 => "0000001100110010",34784 => "0000001100110001",
34785 => "0000001100110001",34786 => "0000001100110001",
34787 => "0000001100110001",34788 => "0000001100110001",
34789 => "0000001100110001",34790 => "0000001100110001",
34791 => "0000001100110001",34792 => "0000001100110001",
34793 => "0000001100110001",34794 => "0000001100110001",
34795 => "0000001100110001",34796 => "0000001100110000",
34797 => "0000001100110000",34798 => "0000001100110000",
34799 => "0000001100110000",34800 => "0000001100110000",
34801 => "0000001100110000",34802 => "0000001100110000",
34803 => "0000001100110000",34804 => "0000001100110000",
34805 => "0000001100110000",34806 => "0000001100110000",
34807 => "0000001100110000",34808 => "0000001100101111",
34809 => "0000001100101111",34810 => "0000001100101111",
34811 => "0000001100101111",34812 => "0000001100101111",
34813 => "0000001100101111",34814 => "0000001100101111",
34815 => "0000001100101111",34816 => "0000000101110000",
34817 => "0000000101001101",34818 => "0000000100101101",
34819 => "0000000100010001",34820 => "0000000011110111",
34821 => "0000000011011111",34822 => "0000000011001010",
34823 => "0000000010110111",34824 => "0000000010100101",
34825 => "0000000000001111",34826 => "0000000101001101",
34827 => "0000000000100001",34828 => "0000000101000110",
34829 => "0000000101000011",34830 => "0000000000100000",
34831 => "0000000100111101",34832 => "0000000100111001",
34833 => "0000000000011111",34834 => "0000000100110011",
34835 => "0000000100110000",34836 => "0000000100101101",
34837 => "0000000100101010",34838 => "0000000100100111",
34839 => "0000000100100100",34840 => "0000000100100001",
34841 => "0000000100011111",34842 => "0000000100011100",
34843 => "0000000100011001",34844 => "0000000100010110",
34845 => "0000000100010011",34846 => "0000000100010001",
34847 => "0000000000011011",34848 => "0000000100001011",
34849 => "0000000100001000",34850 => "0000000100000110",
34851 => "0000000100000011",34852 => "0000000100000001",
34853 => "0000000011111110",34854 => "0000000011111100",
34855 => "0000000011111001",34856 => "0000000011110111",
34857 => "0000000011110100",34858 => "0000000011110010",
34859 => "0000000011101111",34860 => "0000000011101101",
34861 => "0000000011101011",34862 => "0000000011101000",
34863 => "0000000000010111",34864 => "0000000011100100",
34865 => "0000000011100001",34866 => "0000000011011111",
34867 => "0000000011011101",34868 => "0000000011011011",
34869 => "0000000011011001",34870 => "0000000011010110",
34871 => "0000000011010100",34872 => "0000000000010101",
34873 => "0000000011010000",34874 => "0000000011001110",
34875 => "0000000011001100",34876 => "0000000011001010",
34877 => "0000000000000010",34878 => "0000000011000110",
34879 => "0000000011000100",34880 => "0000000011000010",
34881 => "0000000011000000",34882 => "0000000000010011",
34883 => "0000000010111100",34884 => "0000000010111010",
34885 => "0000000010111001",34886 => "0000000010110111",
34887 => "0000000010110101",34888 => "0000000010110011",
34889 => "0000000010110001",34890 => "0000000010110000",
34891 => "0000000010101110",34892 => "0000000010101100",
34893 => "0000000000010001",34894 => "0000000010101001",
34895 => "0000000010100111",34896 => "0000000010100101",
34897 => "0000000010100100",34898 => "0000000010100010",
34899 => "0000000000010000",34900 => "0000000010011111",
34901 => "0000000010011101",34902 => "0000000010011100",
34903 => "0000000010011010",34904 => "0000000010011001",
34905 => "0000000010010111",34906 => "0000000000001111",
34907 => "0000000010010100",34908 => "0000000010010011",
34909 => "0000000010010001",34910 => "0000000010010000",
34911 => "0000000010001110",34912 => "0000000010001101",
34913 => "0000000010001011",34914 => "0000000010001010",
34915 => "0000000010001001",34916 => "0000000101001101",
34917 => "0000000101001101",34918 => "0000000101001100",
34919 => "0000000101001100",34920 => "0000000101001100",
34921 => "0000000101001011",34922 => "0000000101001011",
34923 => "0000000101001011",34924 => "0000000000100001",
34925 => "0000000000100001",34926 => "0000000000100001",
34927 => "0000000101001001",34928 => "0000000101001001",
34929 => "0000000101001001",34930 => "0000000101001000",
34931 => "0000000101001000",34932 => "0000000101001000",
34933 => "0000000101000111",34934 => "0000000101000111",
34935 => "0000000101000111",34936 => "0000000101000110",
34937 => "0000000101000110",34938 => "0000000101000110",
34939 => "0000000101000101",34940 => "0000000101000101",
34941 => "0000000101000101",34942 => "0000000101000100",
34943 => "0000000101000100",34944 => "0000000101000100",
34945 => "0000000101000011",34946 => "0000000101000011",
34947 => "0000000101000011",34948 => "0000000101000010",
34949 => "0000000101000010",34950 => "0000000101000010",
34951 => "0000000101000001",34952 => "0000000101000001",
34953 => "0000000101000001",34954 => "0000000000100000",
34955 => "0000000000100000",34956 => "0000000000100000",
34957 => "0000000100111111",34958 => "0000000100111111",
34959 => "0000000100111111",34960 => "0000000100111111",
34961 => "0000000100111110",34962 => "0000000100111110",
34963 => "0000000100111110",34964 => "0000000100111101",
34965 => "0000000100111101",34966 => "0000000100111101",
34967 => "0000000100111100",34968 => "0000000100111100",
34969 => "0000000100111100",34970 => "0000000100111011",
34971 => "0000000100111011",34972 => "0000000100111011",
34973 => "0000000100111010",34974 => "0000000100111010",
34975 => "0000000100111010",34976 => "0000000100111001",
34977 => "0000000100111001",34978 => "0000000100111001",
34979 => "0000000100111001",34980 => "0000000100111000",
34981 => "0000000100111000",34982 => "0000000100111000",
34983 => "0000000100110111",34984 => "0000000100110111",
34985 => "0000000100110111",34986 => "0000000000011111",
34987 => "0000000000011111",34988 => "0000000000011111",
34989 => "0000000100110101",34990 => "0000000100110101",
34991 => "0000000100110101",34992 => "0000000100110101",
34993 => "0000000100110100",34994 => "0000000100110100",
34995 => "0000000100110100",34996 => "0000000100110011",
34997 => "0000000100110011",34998 => "0000000100110011",
34999 => "0000000100110010",35000 => "0000000100110010",
35001 => "0000000100110010",35002 => "0000000100110001",
35003 => "0000000100110001",35004 => "0000000100110001",
35005 => "0000000100110001",35006 => "0000000100110000",
35007 => "0000000100110000",35008 => "0000000100110000",
35009 => "0000000100101111",35010 => "0000000100101111",
35011 => "0000000100101111",35012 => "0000000100101110",
35013 => "0000000100101110",35014 => "0000000100101110",
35015 => "0000000100101101",35016 => "0000000100101101",
35017 => "0000000100101101",35018 => "0000000100101101",
35019 => "0000000000000011",35020 => "0000000000000011",
35021 => "0000000000000011",35022 => "0000000100101011",
35023 => "0000000100101011",35024 => "0000000100101011",
35025 => "0000000100101010",35026 => "0000000100101010",
35027 => "0000000100101010",35028 => "0000000100101010",
35029 => "0000000100101001",35030 => "0000000100101001",
35031 => "0000000100101001",35032 => "0000000100101000",
35033 => "0000000100101000",35034 => "0000000100101000",
35035 => "0000000100101000",35036 => "0000000100100111",
35037 => "0000000100100111",35038 => "0000000100100111",
35039 => "0000000100100110",35040 => "0000000100100110",
35041 => "0000000100100110",35042 => "0000000100100101",
35043 => "0000000100100101",35044 => "0000000100100101",
35045 => "0000000100100101",35046 => "0000000100100100",
35047 => "0000000100100100",35048 => "0000000100100100",
35049 => "0000000100100011",35050 => "0000000100100011",
35051 => "0000000100100011",35052 => "0000000100100011",
35053 => "0000000000011101",35054 => "0000000000011101",
35055 => "0000000000011101",35056 => "0000000100100001",
35057 => "0000000100100001",35058 => "0000000100100001",
35059 => "0000000100100001",35060 => "0000000100100000",
35061 => "0000000100100000",35062 => "0000000100100000",
35063 => "0000000100011111",35064 => "0000000100011111",
35065 => "0000000100011111",35066 => "0000000100011111",
35067 => "0000000100011110",35068 => "0000000100011110",
35069 => "0000000100011110",35070 => "0000000100011101",
35071 => "0000000100011101",35072 => "0000000100011101",
35073 => "0000000100011101",35074 => "0000000100011100",
35075 => "0000000100011100",35076 => "0000000100011100",
35077 => "0000000100011011",35078 => "0000000100011011",
35079 => "0000000100011011",35080 => "0000000100011011",
35081 => "0000000100011010",35082 => "0000000100011010",
35083 => "0000000100011010",35084 => "0000000100011001",
35085 => "0000000100011001",35086 => "0000000100011001",
35087 => "0000000100011001",35088 => "0000000000011100",
35089 => "0000000000011100",35090 => "0000000000011100",
35091 => "0000000100010111",35092 => "0000000100010111",
35093 => "0000000100010111",35094 => "0000000100010111",
35095 => "0000000100010110",35096 => "0000000100010110",
35097 => "0000000100010110",35098 => "0000000100010101",
35099 => "0000000100010101",35100 => "0000000100010101",
35101 => "0000000100010101",35102 => "0000000100010100",
35103 => "0000000100010100",35104 => "0000000100010100",
35105 => "0000000100010100",35106 => "0000000100010011",
35107 => "0000000100010011",35108 => "0000000100010011",
35109 => "0000000100010010",35110 => "0000000100010010",
35111 => "0000000100010010",35112 => "0000000100010010",
35113 => "0000000100010001",35114 => "0000000100010001",
35115 => "0000000100010001",35116 => "0000000100010001",
35117 => "0000000100010000",35118 => "0000000100010000",
35119 => "0000000100010000",35120 => "0000000100001111",
35121 => "0000000100001111",35122 => "0000000100001111",
35123 => "0000000100001111",35124 => "0000000000011011",
35125 => "0000000000011011",35126 => "0000000000011011",
35127 => "0000000000011011",35128 => "0000000100001101",
35129 => "0000000100001101",35130 => "0000000100001101",
35131 => "0000000100001100",35132 => "0000000100001100",
35133 => "0000000100001100",35134 => "0000000100001100",
35135 => "0000000100001011",35136 => "0000000100001011",
35137 => "0000000100001011",35138 => "0000000100001011",
35139 => "0000000100001010",35140 => "0000000100001010",
35141 => "0000000100001010",35142 => "0000000100001010",
35143 => "0000000100001001",35144 => "0000000100001001",
35145 => "0000000100001001",35146 => "0000000100001000",
35147 => "0000000100001000",35148 => "0000000100001000",
35149 => "0000000100001000",35150 => "0000000100000111",
35151 => "0000000100000111",35152 => "0000000100000111",
35153 => "0000000100000111",35154 => "0000000100000110",
35155 => "0000000100000110",35156 => "0000000100000110",
35157 => "0000000100000110",35158 => "0000000100000101",
35159 => "0000000100000101",35160 => "0000000100000101",
35161 => "0000000100000101",35162 => "0000000000011010",
35163 => "0000000000011010",35164 => "0000000000011010",
35165 => "0000000100000011",35166 => "0000000100000011",
35167 => "0000000100000011",35168 => "0000000100000011",
35169 => "0000000100000010",35170 => "0000000100000010",
35171 => "0000000100000010",35172 => "0000000100000010",
35173 => "0000000100000001",35174 => "0000000100000001",
35175 => "0000000100000001",35176 => "0000000100000001",
35177 => "0000000100000000",35178 => "0000000100000000",
35179 => "0000000100000000",35180 => "0000000100000000",
35181 => "0000000011111111",35182 => "0000000011111111",
35183 => "0000000011111111",35184 => "0000000011111111",
35185 => "0000000011111110",35186 => "0000000011111110",
35187 => "0000000011111110",35188 => "0000000011111110",
35189 => "0000000011111101",35190 => "0000000011111101",
35191 => "0000000011111101",35192 => "0000000011111101",
35193 => "0000000011111100",35194 => "0000000011111100",
35195 => "0000000011111100",35196 => "0000000011111100",
35197 => "0000000011111011",35198 => "0000000011111011",
35199 => "0000000011111011",35200 => "0000000011111011",
35201 => "0000000000011001",35202 => "0000000000011001",
35203 => "0000000000011001",35204 => "0000000000011001",
35205 => "0000000011111001",35206 => "0000000011111001",
35207 => "0000000011111001",35208 => "0000000011111001",
35209 => "0000000011111000",35210 => "0000000011111000",
35211 => "0000000011111000",35212 => "0000000011111000",
35213 => "0000000011110111",35214 => "0000000011110111",
35215 => "0000000011110111",35216 => "0000000011110111",
35217 => "0000000011110110",35218 => "0000000011110110",
35219 => "0000000011110110",35220 => "0000000011110110",
35221 => "0000000011110101",35222 => "0000000011110101",
35223 => "0000000011110101",35224 => "0000000011110101",
35225 => "0000000011110100",35226 => "0000000011110100",
35227 => "0000000011110100",35228 => "0000000011110100",
35229 => "0000000011110011",35230 => "0000000011110011",
35231 => "0000000011110011",35232 => "0000000011110011",
35233 => "0000000011110010",35234 => "0000000011110010",
35235 => "0000000011110010",35236 => "0000000011110010",
35237 => "0000000011110001",35238 => "0000000011110001",
35239 => "0000000011110001",35240 => "0000000011110001",
35241 => "0000000011110001",35242 => "0000000000011000",
35243 => "0000000000011000",35244 => "0000000000011000",
35245 => "0000000000011000",35246 => "0000000011101111",
35247 => "0000000011101111",35248 => "0000000011101111",
35249 => "0000000011101111",35250 => "0000000011101110",
35251 => "0000000011101110",35252 => "0000000011101110",
35253 => "0000000011101110",35254 => "0000000011101101",
35255 => "0000000011101101",35256 => "0000000011101101",
35257 => "0000000011101101",35258 => "0000000011101100",
35259 => "0000000011101100",35260 => "0000000011101100",
35261 => "0000000011101100",35262 => "0000000011101100",
35263 => "0000000011101011",35264 => "0000000011101011",
35265 => "0000000011101011",35266 => "0000000011101011",
35267 => "0000000011101010",35268 => "0000000011101010",
35269 => "0000000011101010",35270 => "0000000011101010",
35271 => "0000000011101001",35272 => "0000000011101001",
35273 => "0000000011101001",35274 => "0000000011101001",
35275 => "0000000011101000",35276 => "0000000011101000",
35277 => "0000000011101000",35278 => "0000000011101000",
35279 => "0000000011101000",35280 => "0000000011100111",
35281 => "0000000011100111",35282 => "0000000011100111",
35283 => "0000000011100111",35284 => "0000000000010111",
35285 => "0000000000010111",35286 => "0000000000010111",
35287 => "0000000000010111",35288 => "0000000011100101",
35289 => "0000000011100101",35290 => "0000000011100101",
35291 => "0000000011100101",35292 => "0000000011100101",
35293 => "0000000011100100",35294 => "0000000011100100",
35295 => "0000000011100100",35296 => "0000000011100100",
35297 => "0000000011100011",35298 => "0000000011100011",
35299 => "0000000011100011",35300 => "0000000011100011",
35301 => "0000000011100011",35302 => "0000000011100010",
35303 => "0000000011100010",35304 => "0000000011100010",
35305 => "0000000011100010",35306 => "0000000011100001",
35307 => "0000000011100001",35308 => "0000000011100001",
35309 => "0000000011100001",35310 => "0000000011100000",
35311 => "0000000011100000",35312 => "0000000011100000",
35313 => "0000000011100000",35314 => "0000000011100000",
35315 => "0000000011011111",35316 => "0000000011011111",
35317 => "0000000011011111",35318 => "0000000011011111",
35319 => "0000000011011110",35320 => "0000000011011110",
35321 => "0000000011011110",35322 => "0000000011011110",
35323 => "0000000011011110",35324 => "0000000011011101",
35325 => "0000000011011101",35326 => "0000000011011101",
35327 => "0000000011011101",35328 => "0000000000010110",
35329 => "0000000000010110",35330 => "0000000000010110",
35331 => "0000000000010110",35332 => "0000000000010110",
35333 => "0000000011011011",35334 => "0000000011011011",
35335 => "0000000011011011",35336 => "0000000011011011",
35337 => "0000000011011010",35338 => "0000000011011010",
35339 => "0000000011011010",35340 => "0000000011011010",
35341 => "0000000011011010",35342 => "0000000011011001",
35343 => "0000000011011001",35344 => "0000000011011001",
35345 => "0000000011011001",35346 => "0000000011011001",
35347 => "0000000011011000",35348 => "0000000011011000",
35349 => "0000000011011000",35350 => "0000000011011000",
35351 => "0000000011010111",35352 => "0000000011010111",
35353 => "0000000011010111",35354 => "0000000011010111",
35355 => "0000000011010111",35356 => "0000000011010110",
35357 => "0000000011010110",35358 => "0000000011010110",
35359 => "0000000011010110",35360 => "0000000011010110",
35361 => "0000000011010101",35362 => "0000000011010101",
35363 => "0000000011010101",35364 => "0000000011010101",
35365 => "0000000011010100",35366 => "0000000011010100",
35367 => "0000000011010100",35368 => "0000000011010100",
35369 => "0000000011010100",35370 => "0000000011010011",
35371 => "0000000011010011",35372 => "0000000011010011",
35373 => "0000000011010011",35374 => "0000000011010011",
35375 => "0000000000010101",35376 => "0000000000010101",
35377 => "0000000000010101",35378 => "0000000000010101",
35379 => "0000000000010101",35380 => "0000000011010001",
35381 => "0000000011010001",35382 => "0000000011010001",
35383 => "0000000011010001",35384 => "0000000011010000",
35385 => "0000000011010000",35386 => "0000000011010000",
35387 => "0000000011010000",35388 => "0000000011010000",
35389 => "0000000011001111",35390 => "0000000011001111",
35391 => "0000000011001111",35392 => "0000000011001111",
35393 => "0000000011001111",35394 => "0000000011001110",
35395 => "0000000011001110",35396 => "0000000011001110",
35397 => "0000000011001110",35398 => "0000000011001110",
35399 => "0000000011001101",35400 => "0000000011001101",
35401 => "0000000011001101",35402 => "0000000011001101",
35403 => "0000000011001101",35404 => "0000000011001100",
35405 => "0000000011001100",35406 => "0000000011001100",
35407 => "0000000011001100",35408 => "0000000011001100",
35409 => "0000000011001011",35410 => "0000000011001011",
35411 => "0000000011001011",35412 => "0000000011001011",
35413 => "0000000011001011",35414 => "0000000011001010",
35415 => "0000000011001010",35416 => "0000000011001010",
35417 => "0000000011001010",35418 => "0000000011001001",
35419 => "0000000011001001",35420 => "0000000011001001",
35421 => "0000000011001001",35422 => "0000000011001001",
35423 => "0000000000000010",35424 => "0000000000000010",
35425 => "0000000000000010",35426 => "0000000000000010",
35427 => "0000000000000010",35428 => "0000000011000111",
35429 => "0000000011000111",35430 => "0000000011000111",
35431 => "0000000011000111",35432 => "0000000011000111",
35433 => "0000000011000110",35434 => "0000000011000110",
35435 => "0000000011000110",35436 => "0000000011000110",
35437 => "0000000011000110",35438 => "0000000011000110",
35439 => "0000000011000101",35440 => "0000000011000101",
35441 => "0000000011000101",35442 => "0000000011000101",
35443 => "0000000011000101",35444 => "0000000011000100",
35445 => "0000000011000100",35446 => "0000000011000100",
35447 => "0000000011000100",35448 => "0000000011000100",
35449 => "0000000011000011",35450 => "0000000011000011",
35451 => "0000000011000011",35452 => "0000000011000011",
35453 => "0000000011000011",35454 => "0000000011000010",
35455 => "0000000011000010",35456 => "0000000011000010",
35457 => "0000000011000010",35458 => "0000000011000010",
35459 => "0000000011000001",35460 => "0000000011000001",
35461 => "0000000011000001",35462 => "0000000011000001",
35463 => "0000000011000001",35464 => "0000000011000000",
35465 => "0000000011000000",35466 => "0000000011000000",
35467 => "0000000011000000",35468 => "0000000011000000",
35469 => "0000000010111111",35470 => "0000000010111111",
35471 => "0000000010111111",35472 => "0000000010111111",
35473 => "0000000010111111",35474 => "0000000010111111",
35475 => "0000000000010011",35476 => "0000000000010011",
35477 => "0000000000010011",35478 => "0000000000010011",
35479 => "0000000000010011",35480 => "0000000010111101",
35481 => "0000000010111101",35482 => "0000000010111101",
35483 => "0000000010111101",35484 => "0000000010111101",
35485 => "0000000010111100",35486 => "0000000010111100",
35487 => "0000000010111100",35488 => "0000000010111100",
35489 => "0000000010111100",35490 => "0000000010111011",
35491 => "0000000010111011",35492 => "0000000010111011",
35493 => "0000000010111011",35494 => "0000000010111011",
35495 => "0000000010111011",35496 => "0000000010111010",
35497 => "0000000010111010",35498 => "0000000010111010",
35499 => "0000000010111010",35500 => "0000000010111010",
35501 => "0000000010111001",35502 => "0000000010111001",
35503 => "0000000010111001",35504 => "0000000010111001",
35505 => "0000000010111001",35506 => "0000000010111001",
35507 => "0000000010111000",35508 => "0000000010111000",
35509 => "0000000010111000",35510 => "0000000010111000",
35511 => "0000000010111000",35512 => "0000000010110111",
35513 => "0000000010110111",35514 => "0000000010110111",
35515 => "0000000010110111",35516 => "0000000010110111",
35517 => "0000000010110111",35518 => "0000000010110110",
35519 => "0000000010110110",35520 => "0000000010110110",
35521 => "0000000010110110",35522 => "0000000010110110",
35523 => "0000000010110101",35524 => "0000000010110101",
35525 => "0000000010110101",35526 => "0000000010110101",
35527 => "0000000010110101",35528 => "0000000010110101",
35529 => "0000000000010010",35530 => "0000000000010010",
35531 => "0000000000010010",35532 => "0000000000010010",
35533 => "0000000000010010",35534 => "0000000010110011",
35535 => "0000000010110011",35536 => "0000000010110011",
35537 => "0000000010110011",35538 => "0000000010110011",
35539 => "0000000010110011",35540 => "0000000010110010",
35541 => "0000000010110010",35542 => "0000000010110010",
35543 => "0000000010110010",35544 => "0000000010110010",
35545 => "0000000010110001",35546 => "0000000010110001",
35547 => "0000000010110001",35548 => "0000000010110001",
35549 => "0000000010110001",35550 => "0000000010110001",
35551 => "0000000010110000",35552 => "0000000010110000",
35553 => "0000000010110000",35554 => "0000000010110000",
35555 => "0000000010110000",35556 => "0000000010110000",
35557 => "0000000010101111",35558 => "0000000010101111",
35559 => "0000000010101111",35560 => "0000000010101111",
35561 => "0000000010101111",35562 => "0000000010101110",
35563 => "0000000010101110",35564 => "0000000010101110",
35565 => "0000000010101110",35566 => "0000000010101110",
35567 => "0000000010101110",35568 => "0000000010101101",
35569 => "0000000010101101",35570 => "0000000010101101",
35571 => "0000000010101101",35572 => "0000000010101101",
35573 => "0000000010101101",35574 => "0000000010101100",
35575 => "0000000010101100",35576 => "0000000010101100",
35577 => "0000000010101100",35578 => "0000000010101100",
35579 => "0000000010101100",35580 => "0000000010101011",
35581 => "0000000010101011",35582 => "0000000010101011",
35583 => "0000000010101011",35584 => "0000000010101011",
35585 => "0000000010101011",35586 => "0000000000010001",
35587 => "0000000000010001",35588 => "0000000000010001",
35589 => "0000000000010001",35590 => "0000000000010001",
35591 => "0000000010101001",35592 => "0000000010101001",
35593 => "0000000010101001",35594 => "0000000010101001",
35595 => "0000000010101001",35596 => "0000000010101001",
35597 => "0000000010101000",35598 => "0000000010101000",
35599 => "0000000010101000",35600 => "0000000010101000",
35601 => "0000000010101000",35602 => "0000000010101000",
35603 => "0000000010100111",35604 => "0000000010100111",
35605 => "0000000010100111",35606 => "0000000010100111",
35607 => "0000000010100111",35608 => "0000000010100111",
35609 => "0000000010100110",35610 => "0000000010100110",
35611 => "0000000010100110",35612 => "0000000010100110",
35613 => "0000000010100110",35614 => "0000000010100110",
35615 => "0000000010100101",35616 => "0000000010100101",
35617 => "0000000010100101",35618 => "0000000010100101",
35619 => "0000000010100101",35620 => "0000000010100101",
35621 => "0000000010100100",35622 => "0000000010100100",
35623 => "0000000010100100",35624 => "0000000010100100",
35625 => "0000000010100100",35626 => "0000000010100100",
35627 => "0000000010100011",35628 => "0000000010100011",
35629 => "0000000010100011",35630 => "0000000010100011",
35631 => "0000000010100011",35632 => "0000000010100011",
35633 => "0000000010100011",35634 => "0000000010100010",
35635 => "0000000010100010",35636 => "0000000010100010",
35637 => "0000000010100010",35638 => "0000000010100010",
35639 => "0000000010100010",35640 => "0000000010100001",
35641 => "0000000010100001",35642 => "0000000010100001",
35643 => "0000000010100001",35644 => "0000000010100001",
35645 => "0000000010100001",35646 => "0000000000010000",
35647 => "0000000000010000",35648 => "0000000000010000",
35649 => "0000000000010000",35650 => "0000000000010000",
35651 => "0000000000010000",35652 => "0000000010011111",
35653 => "0000000010011111",35654 => "0000000010011111",
35655 => "0000000010011111",35656 => "0000000010011111",
35657 => "0000000010011111",35658 => "0000000010011111",
35659 => "0000000010011110",35660 => "0000000010011110",
35661 => "0000000010011110",35662 => "0000000010011110",
35663 => "0000000010011110",35664 => "0000000010011110",
35665 => "0000000010011101",35666 => "0000000010011101",
35667 => "0000000010011101",35668 => "0000000010011101",
35669 => "0000000010011101",35670 => "0000000010011101",
35671 => "0000000010011100",35672 => "0000000010011100",
35673 => "0000000010011100",35674 => "0000000010011100",
35675 => "0000000010011100",35676 => "0000000010011100",
35677 => "0000000010011100",35678 => "0000000010011011",
35679 => "0000000010011011",35680 => "0000000010011011",
35681 => "0000000010011011",35682 => "0000000010011011",
35683 => "0000000010011011",35684 => "0000000010011010",
35685 => "0000000010011010",35686 => "0000000010011010",
35687 => "0000000010011010",35688 => "0000000010011010",
35689 => "0000000010011010",35690 => "0000000010011010",
35691 => "0000000010011001",35692 => "0000000010011001",
35693 => "0000000010011001",35694 => "0000000010011001",
35695 => "0000000010011001",35696 => "0000000010011001",
35697 => "0000000010011000",35698 => "0000000010011000",
35699 => "0000000010011000",35700 => "0000000010011000",
35701 => "0000000010011000",35702 => "0000000010011000",
35703 => "0000000010011000",35704 => "0000000010010111",
35705 => "0000000010010111",35706 => "0000000010010111",
35707 => "0000000010010111",35708 => "0000000010010111",
35709 => "0000000010010111",35710 => "0000000000001111",
35711 => "0000000000001111",35712 => "0000000000001111",
35713 => "0000000000001111",35714 => "0000000000001111",
35715 => "0000000000001111",35716 => "0000000000001111",
35717 => "0000000010010101",35718 => "0000000010010101",
35719 => "0000000010010101",35720 => "0000000010010101",
35721 => "0000000010010101",35722 => "0000000010010101",
35723 => "0000000010010101",35724 => "0000000010010100",
35725 => "0000000010010100",35726 => "0000000010010100",
35727 => "0000000010010100",35728 => "0000000010010100",
35729 => "0000000010010100",35730 => "0000000010010011",
35731 => "0000000010010011",35732 => "0000000010010011",
35733 => "0000000010010011",35734 => "0000000010010011",
35735 => "0000000010010011",35736 => "0000000010010011",
35737 => "0000000010010010",35738 => "0000000010010010",
35739 => "0000000010010010",35740 => "0000000010010010",
35741 => "0000000010010010",35742 => "0000000010010010",
35743 => "0000000010010010",35744 => "0000000010010001",
35745 => "0000000010010001",35746 => "0000000010010001",
35747 => "0000000010010001",35748 => "0000000010010001",
35749 => "0000000010010001",35750 => "0000000010010001",
35751 => "0000000010010000",35752 => "0000000010010000",
35753 => "0000000010010000",35754 => "0000000010010000",
35755 => "0000000010010000",35756 => "0000000010010000",
35757 => "0000000010010000",35758 => "0000000010001111",
35759 => "0000000010001111",35760 => "0000000010001111",
35761 => "0000000010001111",35762 => "0000000010001111",
35763 => "0000000010001111",35764 => "0000000010001111",
35765 => "0000000010001110",35766 => "0000000010001110",
35767 => "0000000010001110",35768 => "0000000010001110",
35769 => "0000000010001110",35770 => "0000000010001110",
35771 => "0000000010001110",35772 => "0000000010001101",
35773 => "0000000010001101",35774 => "0000000010001101",
35775 => "0000000010001101",35776 => "0000000010001101",
35777 => "0000000010001101",35778 => "0000000010001101",
35779 => "0000000000001110",35780 => "0000000000001110",
35781 => "0000000000001110",35782 => "0000000000001110",
35783 => "0000000000001110",35784 => "0000000000001110",
35785 => "0000000000001110",35786 => "0000000010001011",
35787 => "0000000010001011",35788 => "0000000010001011",
35789 => "0000000010001011",35790 => "0000000010001011",
35791 => "0000000010001011",35792 => "0000000010001011",
35793 => "0000000010001010",35794 => "0000000010001010",
35795 => "0000000010001010",35796 => "0000000010001010",
35797 => "0000000010001010",35798 => "0000000010001010",
35799 => "0000000010001010",35800 => "0000000010001010",
35801 => "0000000010001001",35802 => "0000000010001001",
35803 => "0000000010001001",35804 => "0000000010001001",
35805 => "0000000010001001",35806 => "0000000010001001",
35807 => "0000000010001001",35808 => "0000000010001000",
35809 => "0000000010001000",35810 => "0000000010001000",
35811 => "0000000010001000",35812 => "0000000010001000",
35813 => "0000000010001000",35814 => "0000000010001000",
35815 => "0000000010000111",35816 => "0000000101001101",
35817 => "0000000101001101",35818 => "0000000101001101",
35819 => "0000000101001101",35820 => "0000000101001101",
35821 => "0000000101001101",35822 => "0000000101001101",
35823 => "0000000101001101",35824 => "0000000101001101",
35825 => "0000000101001101",35826 => "0000000101001101",
35827 => "0000000101001101",35828 => "0000000101001100",
35829 => "0000000101001100",35830 => "0000000101001100",
35831 => "0000000101001100",35832 => "0000000101001100",
35833 => "0000000101001100",35834 => "0000000101001100",
35835 => "0000000101001100",35836 => "0000000101001100",
35837 => "0000000101001100",35838 => "0000000101001100",
35839 => "0000000101001100",35840 => "0000000101001100",
35841 => "0000000101001100",35842 => "0000000101001100",
35843 => "0000000101001100",35844 => "0000000101001100",
35845 => "0000000101001100",35846 => "0000000101001100",
35847 => "0000000101001100",35848 => "0000000101001100",
35849 => "0000000101001100",35850 => "0000000101001100",
35851 => "0000000101001100",35852 => "0000000101001100",
35853 => "0000000101001100",35854 => "0000000101001100",
35855 => "0000000101001100",35856 => "0000000101001100",
35857 => "0000000101001100",35858 => "0000000101001011",
35859 => "0000000101001011",35860 => "0000000101001011",
35861 => "0000000101001011",35862 => "0000000101001011",
35863 => "0000000101001011",35864 => "0000000101001011",
35865 => "0000000101001011",35866 => "0000000101001011",
35867 => "0000000101001011",35868 => "0000000101001011",
35869 => "0000000101001011",35870 => "0000000101001011",
35871 => "0000000101001011",35872 => "0000000101001011",
35873 => "0000000101001011",35874 => "0000000101001011",
35875 => "0000000101001011",35876 => "0000000101001011",
35877 => "0000000101001011",35878 => "0000000101001011",
35879 => "0000000101001011",35880 => "0000000101001011",
35881 => "0000000101001011",35882 => "0000000101001011",
35883 => "0000000101001011",35884 => "0000000101001011",
35885 => "0000000101001011",35886 => "0000000101001011",
35887 => "0000000101001011",35888 => "0000000000100001",
35889 => "0000000000100001",35890 => "0000000000100001",
35891 => "0000000000100001",35892 => "0000000000100001",
35893 => "0000000000100001",35894 => "0000000000100001",
35895 => "0000000000100001",35896 => "0000000000100001",
35897 => "0000000000100001",35898 => "0000000000100001",
35899 => "0000000000100001",35900 => "0000000000100001",
35901 => "0000000000100001",35902 => "0000000000100001",
35903 => "0000000000100001",35904 => "0000000000100001",
35905 => "0000000000100001",35906 => "0000000000100001",
35907 => "0000000000100001",35908 => "0000000000100001",
35909 => "0000000000100001",35910 => "0000000000100001",
35911 => "0000000000100001",35912 => "0000000000100001",
35913 => "0000000000100001",35914 => "0000000000100001",
35915 => "0000000000100001",35916 => "0000000000100001",
35917 => "0000000000100001",35918 => "0000000101001001",
35919 => "0000000101001001",35920 => "0000000101001001",
35921 => "0000000101001001",35922 => "0000000101001001",
35923 => "0000000101001001",35924 => "0000000101001001",
35925 => "0000000101001001",35926 => "0000000101001001",
35927 => "0000000101001001",35928 => "0000000101001001",
35929 => "0000000101001001",35930 => "0000000101001001",
35931 => "0000000101001001",35932 => "0000000101001001",
35933 => "0000000101001001",35934 => "0000000101001001",
35935 => "0000000101001001",35936 => "0000000101001001",
35937 => "0000000101001001",35938 => "0000000101001001",
35939 => "0000000101001001",35940 => "0000000101001001",
35941 => "0000000101001001",35942 => "0000000101001001",
35943 => "0000000101001001",35944 => "0000000101001001",
35945 => "0000000101001001",35946 => "0000000101001001",
35947 => "0000000101001001",35948 => "0000000101001001",
35949 => "0000000101001000",35950 => "0000000101001000",
35951 => "0000000101001000",35952 => "0000000101001000",
35953 => "0000000101001000",35954 => "0000000101001000",
35955 => "0000000101001000",35956 => "0000000101001000",
35957 => "0000000101001000",35958 => "0000000101001000",
35959 => "0000000101001000",35960 => "0000000101001000",
35961 => "0000000101001000",35962 => "0000000101001000",
35963 => "0000000101001000",35964 => "0000000101001000",
35965 => "0000000101001000",35966 => "0000000101001000",
35967 => "0000000101001000",35968 => "0000000101001000",
35969 => "0000000101001000",35970 => "0000000101001000",
35971 => "0000000101001000",35972 => "0000000101001000",
35973 => "0000000101001000",35974 => "0000000101001000",
35975 => "0000000101001000",35976 => "0000000101001000",
35977 => "0000000101001000",35978 => "0000000101001000",
35979 => "0000000101000111",35980 => "0000000101000111",
35981 => "0000000101000111",35982 => "0000000101000111",
35983 => "0000000101000111",35984 => "0000000101000111",
35985 => "0000000101000111",35986 => "0000000101000111",
35987 => "0000000101000111",35988 => "0000000101000111",
35989 => "0000000101000111",35990 => "0000000101000111",
35991 => "0000000101000111",35992 => "0000000101000111",
35993 => "0000000101000111",35994 => "0000000101000111",
35995 => "0000000101000111",35996 => "0000000101000111",
35997 => "0000000101000111",35998 => "0000000101000111",
35999 => "0000000101000111",36000 => "0000000101000111",
36001 => "0000000101000111",36002 => "0000000101000111",
36003 => "0000000101000111",36004 => "0000000101000111",
36005 => "0000000101000111",36006 => "0000000101000111",
36007 => "0000000101000111",36008 => "0000000101000111",
36009 => "0000000101000111",36010 => "0000000101000110",
36011 => "0000000101000110",36012 => "0000000101000110",
36013 => "0000000101000110",36014 => "0000000101000110",
36015 => "0000000101000110",36016 => "0000000101000110",
36017 => "0000000101000110",36018 => "0000000101000110",
36019 => "0000000101000110",36020 => "0000000101000110",
36021 => "0000000101000110",36022 => "0000000101000110",
36023 => "0000000101000110",36024 => "0000000101000110",
36025 => "0000000101000110",36026 => "0000000101000110",
36027 => "0000000101000110",36028 => "0000000101000110",
36029 => "0000000101000110",36030 => "0000000101000110",
36031 => "0000000101000110",36032 => "0000000101000110",
36033 => "0000000101000110",36034 => "0000000101000110",
36035 => "0000000101000110",36036 => "0000000101000110",
36037 => "0000000101000110",36038 => "0000000101000110",
36039 => "0000000101000110",36040 => "0000000101000101",
36041 => "0000000101000101",36042 => "0000000101000101",
36043 => "0000000101000101",36044 => "0000000101000101",
36045 => "0000000101000101",36046 => "0000000101000101",
36047 => "0000000101000101",36048 => "0000000101000101",
36049 => "0000000101000101",36050 => "0000000101000101",
36051 => "0000000101000101",36052 => "0000000101000101",
36053 => "0000000101000101",36054 => "0000000101000101",
36055 => "0000000101000101",36056 => "0000000101000101",
36057 => "0000000101000101",36058 => "0000000101000101",
36059 => "0000000101000101",36060 => "0000000101000101",
36061 => "0000000101000101",36062 => "0000000101000101",
36063 => "0000000101000101",36064 => "0000000101000101",
36065 => "0000000101000101",36066 => "0000000101000101",
36067 => "0000000101000101",36068 => "0000000101000101",
36069 => "0000000101000101",36070 => "0000000101000101",
36071 => "0000000101000100",36072 => "0000000101000100",
36073 => "0000000101000100",36074 => "0000000101000100",
36075 => "0000000101000100",36076 => "0000000101000100",
36077 => "0000000101000100",36078 => "0000000101000100",
36079 => "0000000101000100",36080 => "0000000101000100",
36081 => "0000000101000100",36082 => "0000000101000100",
36083 => "0000000101000100",36084 => "0000000101000100",
36085 => "0000000101000100",36086 => "0000000101000100",
36087 => "0000000101000100",36088 => "0000000101000100",
36089 => "0000000101000100",36090 => "0000000101000100",
36091 => "0000000101000100",36092 => "0000000101000100",
36093 => "0000000101000100",36094 => "0000000101000100",
36095 => "0000000101000100",36096 => "0000000101000100",
36097 => "0000000101000100",36098 => "0000000101000100",
36099 => "0000000101000100",36100 => "0000000101000100",
36101 => "0000000101000100",36102 => "0000000101000011",
36103 => "0000000101000011",36104 => "0000000101000011",
36105 => "0000000101000011",36106 => "0000000101000011",
36107 => "0000000101000011",36108 => "0000000101000011",
36109 => "0000000101000011",36110 => "0000000101000011",
36111 => "0000000101000011",36112 => "0000000101000011",
36113 => "0000000101000011",36114 => "0000000101000011",
36115 => "0000000101000011",36116 => "0000000101000011",
36117 => "0000000101000011",36118 => "0000000101000011",
36119 => "0000000101000011",36120 => "0000000101000011",
36121 => "0000000101000011",36122 => "0000000101000011",
36123 => "0000000101000011",36124 => "0000000101000011",
36125 => "0000000101000011",36126 => "0000000101000011",
36127 => "0000000101000011",36128 => "0000000101000011",
36129 => "0000000101000011",36130 => "0000000101000011",
36131 => "0000000101000011",36132 => "0000000101000011",
36133 => "0000000101000010",36134 => "0000000101000010",
36135 => "0000000101000010",36136 => "0000000101000010",
36137 => "0000000101000010",36138 => "0000000101000010",
36139 => "0000000101000010",36140 => "0000000101000010",
36141 => "0000000101000010",36142 => "0000000101000010",
36143 => "0000000101000010",36144 => "0000000101000010",
36145 => "0000000101000010",36146 => "0000000101000010",
36147 => "0000000101000010",36148 => "0000000101000010",
36149 => "0000000101000010",36150 => "0000000101000010",
36151 => "0000000101000010",36152 => "0000000101000010",
36153 => "0000000101000010",36154 => "0000000101000010",
36155 => "0000000101000010",36156 => "0000000101000010",
36157 => "0000000101000010",36158 => "0000000101000010",
36159 => "0000000101000010",36160 => "0000000101000010",
36161 => "0000000101000010",36162 => "0000000101000010",
36163 => "0000000101000010",36164 => "0000000101000001",
36165 => "0000000101000001",36166 => "0000000101000001",
36167 => "0000000101000001",36168 => "0000000101000001",
36169 => "0000000101000001",36170 => "0000000101000001",
36171 => "0000000101000001",36172 => "0000000101000001",
36173 => "0000000101000001",36174 => "0000000101000001",
36175 => "0000000101000001",36176 => "0000000101000001",
36177 => "0000000101000001",36178 => "0000000101000001",
36179 => "0000000101000001",36180 => "0000000101000001",
36181 => "0000000101000001",36182 => "0000000101000001",
36183 => "0000000101000001",36184 => "0000000101000001",
36185 => "0000000101000001",36186 => "0000000101000001",
36187 => "0000000101000001",36188 => "0000000101000001",
36189 => "0000000101000001",36190 => "0000000101000001",
36191 => "0000000101000001",36192 => "0000000101000001",
36193 => "0000000101000001",36194 => "0000000101000001",
36195 => "0000000000100000",36196 => "0000000000100000",
36197 => "0000000000100000",36198 => "0000000000100000",
36199 => "0000000000100000",36200 => "0000000000100000",
36201 => "0000000000100000",36202 => "0000000000100000",
36203 => "0000000000100000",36204 => "0000000000100000",
36205 => "0000000000100000",36206 => "0000000000100000",
36207 => "0000000000100000",36208 => "0000000000100000",
36209 => "0000000000100000",36210 => "0000000000100000",
36211 => "0000000000100000",36212 => "0000000000100000",
36213 => "0000000000100000",36214 => "0000000000100000",
36215 => "0000000000100000",36216 => "0000000000100000",
36217 => "0000000000100000",36218 => "0000000000100000",
36219 => "0000000000100000",36220 => "0000000000100000",
36221 => "0000000000100000",36222 => "0000000000100000",
36223 => "0000000000100000",36224 => "0000000000100000",
36225 => "0000000000100000",36226 => "0000000100111111",
36227 => "0000000100111111",36228 => "0000000100111111",
36229 => "0000000100111111",36230 => "0000000100111111",
36231 => "0000000100111111",36232 => "0000000100111111",
36233 => "0000000100111111",36234 => "0000000100111111",
36235 => "0000000100111111",36236 => "0000000100111111",
36237 => "0000000100111111",36238 => "0000000100111111",
36239 => "0000000100111111",36240 => "0000000100111111",
36241 => "0000000100111111",36242 => "0000000100111111",
36243 => "0000000100111111",36244 => "0000000100111111",
36245 => "0000000100111111",36246 => "0000000100111111",
36247 => "0000000100111111",36248 => "0000000100111111",
36249 => "0000000100111111",36250 => "0000000100111111",
36251 => "0000000100111111",36252 => "0000000100111111",
36253 => "0000000100111111",36254 => "0000000100111111",
36255 => "0000000100111111",36256 => "0000000100111111",
36257 => "0000000100111111",36258 => "0000000100111110",
36259 => "0000000100111110",36260 => "0000000100111110",
36261 => "0000000100111110",36262 => "0000000100111110",
36263 => "0000000100111110",36264 => "0000000100111110",
36265 => "0000000100111110",36266 => "0000000100111110",
36267 => "0000000100111110",36268 => "0000000100111110",
36269 => "0000000100111110",36270 => "0000000100111110",
36271 => "0000000100111110",36272 => "0000000100111110",
36273 => "0000000100111110",36274 => "0000000100111110",
36275 => "0000000100111110",36276 => "0000000100111110",
36277 => "0000000100111110",36278 => "0000000100111110",
36279 => "0000000100111110",36280 => "0000000100111110",
36281 => "0000000100111110",36282 => "0000000100111110",
36283 => "0000000100111110",36284 => "0000000100111110",
36285 => "0000000100111110",36286 => "0000000100111110",
36287 => "0000000100111110",36288 => "0000000100111110",
36289 => "0000000100111101",36290 => "0000000100111101",
36291 => "0000000100111101",36292 => "0000000100111101",
36293 => "0000000100111101",36294 => "0000000100111101",
36295 => "0000000100111101",36296 => "0000000100111101",
36297 => "0000000100111101",36298 => "0000000100111101",
36299 => "0000000100111101",36300 => "0000000100111101",
36301 => "0000000100111101",36302 => "0000000100111101",
36303 => "0000000100111101",36304 => "0000000100111101",
36305 => "0000000100111101",36306 => "0000000100111101",
36307 => "0000000100111101",36308 => "0000000100111101",
36309 => "0000000100111101",36310 => "0000000100111101",
36311 => "0000000100111101",36312 => "0000000100111101",
36313 => "0000000100111101",36314 => "0000000100111101",
36315 => "0000000100111101",36316 => "0000000100111101",
36317 => "0000000100111101",36318 => "0000000100111101",
36319 => "0000000100111101",36320 => "0000000100111101",
36321 => "0000000100111100",36322 => "0000000100111100",
36323 => "0000000100111100",36324 => "0000000100111100",
36325 => "0000000100111100",36326 => "0000000100111100",
36327 => "0000000100111100",36328 => "0000000100111100",
36329 => "0000000100111100",36330 => "0000000100111100",
36331 => "0000000100111100",36332 => "0000000100111100",
36333 => "0000000100111100",36334 => "0000000100111100",
36335 => "0000000100111100",36336 => "0000000100111100",
36337 => "0000000100111100",36338 => "0000000100111100",
36339 => "0000000100111100",36340 => "0000000100111100",
36341 => "0000000100111100",36342 => "0000000100111100",
36343 => "0000000100111100",36344 => "0000000100111100",
36345 => "0000000100111100",36346 => "0000000100111100",
36347 => "0000000100111100",36348 => "0000000100111100",
36349 => "0000000100111100",36350 => "0000000100111100",
36351 => "0000000100111100",36352 => "0000000100111011",
36353 => "0000000100111011",36354 => "0000000100111011",
36355 => "0000000100111011",36356 => "0000000100111011",
36357 => "0000000100111011",36358 => "0000000100111011",
36359 => "0000000100111011",36360 => "0000000100111011",
36361 => "0000000100111011",36362 => "0000000100111011",
36363 => "0000000100111011",36364 => "0000000100111011",
36365 => "0000000100111011",36366 => "0000000100111011",
36367 => "0000000100111011",36368 => "0000000100111011",
36369 => "0000000100111011",36370 => "0000000100111011",
36371 => "0000000100111011",36372 => "0000000100111011",
36373 => "0000000100111011",36374 => "0000000100111011",
36375 => "0000000100111011",36376 => "0000000100111011",
36377 => "0000000100111011",36378 => "0000000100111011",
36379 => "0000000100111011",36380 => "0000000100111011",
36381 => "0000000100111011",36382 => "0000000100111011",
36383 => "0000000100111011",36384 => "0000000100111010",
36385 => "0000000100111010",36386 => "0000000100111010",
36387 => "0000000100111010",36388 => "0000000100111010",
36389 => "0000000100111010",36390 => "0000000100111010",
36391 => "0000000100111010",36392 => "0000000100111010",
36393 => "0000000100111010",36394 => "0000000100111010",
36395 => "0000000100111010",36396 => "0000000100111010",
36397 => "0000000100111010",36398 => "0000000100111010",
36399 => "0000000100111010",36400 => "0000000100111010",
36401 => "0000000100111010",36402 => "0000000100111010",
36403 => "0000000100111010",36404 => "0000000100111010",
36405 => "0000000100111010",36406 => "0000000100111010",
36407 => "0000000100111010",36408 => "0000000100111010",
36409 => "0000000100111010",36410 => "0000000100111010",
36411 => "0000000100111010",36412 => "0000000100111010",
36413 => "0000000100111010",36414 => "0000000100111010",
36415 => "0000000100111010",36416 => "0000000100111001",
36417 => "0000000100111001",36418 => "0000000100111001",
36419 => "0000000100111001",36420 => "0000000100111001",
36421 => "0000000100111001",36422 => "0000000100111001",
36423 => "0000000100111001",36424 => "0000000100111001",
36425 => "0000000100111001",36426 => "0000000100111001",
36427 => "0000000100111001",36428 => "0000000100111001",
36429 => "0000000100111001",36430 => "0000000100111001",
36431 => "0000000100111001",36432 => "0000000100111001",
36433 => "0000000100111001",36434 => "0000000100111001",
36435 => "0000000100111001",36436 => "0000000100111001",
36437 => "0000000100111001",36438 => "0000000100111001",
36439 => "0000000100111001",36440 => "0000000100111001",
36441 => "0000000100111001",36442 => "0000000100111001",
36443 => "0000000100111001",36444 => "0000000100111001",
36445 => "0000000100111001",36446 => "0000000100111001",
36447 => "0000000100111001",36448 => "0000000100111000",
36449 => "0000000100111000",36450 => "0000000100111000",
36451 => "0000000100111000",36452 => "0000000100111000",
36453 => "0000000100111000",36454 => "0000000100111000",
36455 => "0000000100111000",36456 => "0000000100111000",
36457 => "0000000100111000",36458 => "0000000100111000",
36459 => "0000000100111000",36460 => "0000000100111000",
36461 => "0000000100111000",36462 => "0000000100111000",
36463 => "0000000100111000",36464 => "0000000100111000",
36465 => "0000000100111000",36466 => "0000000100111000",
36467 => "0000000100111000",36468 => "0000000100111000",
36469 => "0000000100111000",36470 => "0000000100111000",
36471 => "0000000100111000",36472 => "0000000100111000",
36473 => "0000000100111000",36474 => "0000000100111000",
36475 => "0000000100111000",36476 => "0000000100111000",
36477 => "0000000100111000",36478 => "0000000100111000",
36479 => "0000000100111000",36480 => "0000000100110111",
36481 => "0000000100110111",36482 => "0000000100110111",
36483 => "0000000100110111",36484 => "0000000100110111",
36485 => "0000000100110111",36486 => "0000000100110111",
36487 => "0000000100110111",36488 => "0000000100110111",
36489 => "0000000100110111",36490 => "0000000100110111",
36491 => "0000000100110111",36492 => "0000000100110111",
36493 => "0000000100110111",36494 => "0000000100110111",
36495 => "0000000100110111",36496 => "0000000100110111",
36497 => "0000000100110111",36498 => "0000000100110111",
36499 => "0000000100110111",36500 => "0000000100110111",
36501 => "0000000100110111",36502 => "0000000100110111",
36503 => "0000000100110111",36504 => "0000000100110111",
36505 => "0000000100110111",36506 => "0000000100110111",
36507 => "0000000100110111",36508 => "0000000100110111",
36509 => "0000000100110111",36510 => "0000000100110111",
36511 => "0000000100110111",36512 => "0000000000011111",
36513 => "0000000000011111",36514 => "0000000000011111",
36515 => "0000000000011111",36516 => "0000000000011111",
36517 => "0000000000011111",36518 => "0000000000011111",
36519 => "0000000000011111",36520 => "0000000000011111",
36521 => "0000000000011111",36522 => "0000000000011111",
36523 => "0000000000011111",36524 => "0000000000011111",
36525 => "0000000000011111",36526 => "0000000000011111",
36527 => "0000000000011111",36528 => "0000000000011111",
36529 => "0000000000011111",36530 => "0000000000011111",
36531 => "0000000000011111",36532 => "0000000000011111",
36533 => "0000000000011111",36534 => "0000000000011111",
36535 => "0000000000011111",36536 => "0000000000011111",
36537 => "0000000000011111",36538 => "0000000000011111",
36539 => "0000000000011111",36540 => "0000000000011111",
36541 => "0000000000011111",36542 => "0000000000011111",
36543 => "0000000000011111",36544 => "0000000100110101",
36545 => "0000000100110101",36546 => "0000000100110101",
36547 => "0000000100110101",36548 => "0000000100110101",
36549 => "0000000100110101",36550 => "0000000100110101",
36551 => "0000000100110101",36552 => "0000000100110101",
36553 => "0000000100110101",36554 => "0000000100110101",
36555 => "0000000100110101",36556 => "0000000100110101",
36557 => "0000000100110101",36558 => "0000000100110101",
36559 => "0000000100110101",36560 => "0000000100110101",
36561 => "0000000100110101",36562 => "0000000100110101",
36563 => "0000000100110101",36564 => "0000000100110101",
36565 => "0000000100110101",36566 => "0000000100110101",
36567 => "0000000100110101",36568 => "0000000100110101",
36569 => "0000000100110101",36570 => "0000000100110101",
36571 => "0000000100110101",36572 => "0000000100110101",
36573 => "0000000100110101",36574 => "0000000100110101",
36575 => "0000000100110101",36576 => "0000000100110101",
36577 => "0000000100110100",36578 => "0000000100110100",
36579 => "0000000100110100",36580 => "0000000100110100",
36581 => "0000000100110100",36582 => "0000000100110100",
36583 => "0000000100110100",36584 => "0000000100110100",
36585 => "0000000100110100",36586 => "0000000100110100",
36587 => "0000000100110100",36588 => "0000000100110100",
36589 => "0000000100110100",36590 => "0000000100110100",
36591 => "0000000100110100",36592 => "0000000100110100",
36593 => "0000000100110100",36594 => "0000000100110100",
36595 => "0000000100110100",36596 => "0000000100110100",
36597 => "0000000100110100",36598 => "0000000100110100",
36599 => "0000000100110100",36600 => "0000000100110100",
36601 => "0000000100110100",36602 => "0000000100110100",
36603 => "0000000100110100",36604 => "0000000100110100",
36605 => "0000000100110100",36606 => "0000000100110100",
36607 => "0000000100110100",36608 => "0000000100110100",
36609 => "0000000100110011",36610 => "0000000100110011",
36611 => "0000000100110011",36612 => "0000000100110011",
36613 => "0000000100110011",36614 => "0000000100110011",
36615 => "0000000100110011",36616 => "0000000100110011",
36617 => "0000000100110011",36618 => "0000000100110011",
36619 => "0000000100110011",36620 => "0000000100110011",
36621 => "0000000100110011",36622 => "0000000100110011",
36623 => "0000000100110011",36624 => "0000000100110011",
36625 => "0000000100110011",36626 => "0000000100110011",
36627 => "0000000100110011",36628 => "0000000100110011",
36629 => "0000000100110011",36630 => "0000000100110011",
36631 => "0000000100110011",36632 => "0000000100110011",
36633 => "0000000100110011",36634 => "0000000100110011",
36635 => "0000000100110011",36636 => "0000000100110011",
36637 => "0000000100110011",36638 => "0000000100110011",
36639 => "0000000100110011",36640 => "0000000100110011",
36641 => "0000000100110011",36642 => "0000000100110010",
36643 => "0000000100110010",36644 => "0000000100110010",
36645 => "0000000100110010",36646 => "0000000100110010",
36647 => "0000000100110010",36648 => "0000000100110010",
36649 => "0000000100110010",36650 => "0000000100110010",
36651 => "0000000100110010",36652 => "0000000100110010",
36653 => "0000000100110010",36654 => "0000000100110010",
36655 => "0000000100110010",36656 => "0000000100110010",
36657 => "0000000100110010",36658 => "0000000100110010",
36659 => "0000000100110010",36660 => "0000000100110010",
36661 => "0000000100110010",36662 => "0000000100110010",
36663 => "0000000100110010",36664 => "0000000100110010",
36665 => "0000000100110010",36666 => "0000000100110010",
36667 => "0000000100110010",36668 => "0000000100110010",
36669 => "0000000100110010",36670 => "0000000100110010",
36671 => "0000000100110010",36672 => "0000000100110010",
36673 => "0000000100110010",36674 => "0000000100110010",
36675 => "0000000100110001",36676 => "0000000100110001",
36677 => "0000000100110001",36678 => "0000000100110001",
36679 => "0000000100110001",36680 => "0000000100110001",
36681 => "0000000100110001",36682 => "0000000100110001",
36683 => "0000000100110001",36684 => "0000000100110001",
36685 => "0000000100110001",36686 => "0000000100110001",
36687 => "0000000100110001",36688 => "0000000100110001",
36689 => "0000000100110001",36690 => "0000000100110001",
36691 => "0000000100110001",36692 => "0000000100110001",
36693 => "0000000100110001",36694 => "0000000100110001",
36695 => "0000000100110001",36696 => "0000000100110001",
36697 => "0000000100110001",36698 => "0000000100110001",
36699 => "0000000100110001",36700 => "0000000100110001",
36701 => "0000000100110001",36702 => "0000000100110001",
36703 => "0000000100110001",36704 => "0000000100110001",
36705 => "0000000100110001",36706 => "0000000100110001",
36707 => "0000000100110000",36708 => "0000000100110000",
36709 => "0000000100110000",36710 => "0000000100110000",
36711 => "0000000100110000",36712 => "0000000100110000",
36713 => "0000000100110000",36714 => "0000000100110000",
36715 => "0000000100110000",36716 => "0000000100110000",
36717 => "0000000100110000",36718 => "0000000100110000",
36719 => "0000000100110000",36720 => "0000000100110000",
36721 => "0000000100110000",36722 => "0000000100110000",
36723 => "0000000100110000",36724 => "0000000100110000",
36725 => "0000000100110000",36726 => "0000000100110000",
36727 => "0000000100110000",36728 => "0000000100110000",
36729 => "0000000100110000",36730 => "0000000100110000",
36731 => "0000000100110000",36732 => "0000000100110000",
36733 => "0000000100110000",36734 => "0000000100110000",
36735 => "0000000100110000",36736 => "0000000100110000",
36737 => "0000000100110000",36738 => "0000000100110000",
36739 => "0000000100110000",36740 => "0000000100101111",
36741 => "0000000100101111",36742 => "0000000100101111",
36743 => "0000000100101111",36744 => "0000000100101111",
36745 => "0000000100101111",36746 => "0000000100101111",
36747 => "0000000100101111",36748 => "0000000100101111",
36749 => "0000000100101111",36750 => "0000000100101111",
36751 => "0000000100101111",36752 => "0000000100101111",
36753 => "0000000100101111",36754 => "0000000100101111",
36755 => "0000000100101111",36756 => "0000000100101111",
36757 => "0000000100101111",36758 => "0000000100101111",
36759 => "0000000100101111",36760 => "0000000100101111",
36761 => "0000000100101111",36762 => "0000000100101111",
36763 => "0000000100101111",36764 => "0000000100101111",
36765 => "0000000100101111",36766 => "0000000100101111",
36767 => "0000000100101111",36768 => "0000000100101111",
36769 => "0000000100101111",36770 => "0000000100101111",
36771 => "0000000100101111",36772 => "0000000100101111",
36773 => "0000000100101110",36774 => "0000000100101110",
36775 => "0000000100101110",36776 => "0000000100101110",
36777 => "0000000100101110",36778 => "0000000100101110",
36779 => "0000000100101110",36780 => "0000000100101110",
36781 => "0000000100101110",36782 => "0000000100101110",
36783 => "0000000100101110",36784 => "0000000100101110",
36785 => "0000000100101110",36786 => "0000000100101110",
36787 => "0000000100101110",36788 => "0000000100101110",
36789 => "0000000100101110",36790 => "0000000100101110",
36791 => "0000000100101110",36792 => "0000000100101110",
36793 => "0000000100101110",36794 => "0000000100101110",
36795 => "0000000100101110",36796 => "0000000100101110",
36797 => "0000000100101110",36798 => "0000000100101110",
36799 => "0000000100101110",36800 => "0000000100101110",
36801 => "0000000100101110",36802 => "0000000100101110",
36803 => "0000000100101110",36804 => "0000000100101110",
36805 => "0000000100101110",36806 => "0000000100101101",
36807 => "0000000100101101",36808 => "0000000100101101",
36809 => "0000000100101101",36810 => "0000000100101101",
36811 => "0000000100101101",36812 => "0000000100101101",
36813 => "0000000100101101",36814 => "0000000100101101",
36815 => "0000000100101101",36816 => "0000000100101101",
36817 => "0000000100101101",36818 => "0000000100101101",
36819 => "0000000100101101",36820 => "0000000100101101",
36821 => "0000000100101101",36822 => "0000000100101101",
36823 => "0000000100101101",36824 => "0000000100101101",
36825 => "0000000100101101",36826 => "0000000100101101",
36827 => "0000000100101101",36828 => "0000000100101101",
36829 => "0000000100101101",36830 => "0000000100101101",
36831 => "0000000100101101",36832 => "0000000100101101",
36833 => "0000000100101101",36834 => "0000000100101101",
36835 => "0000000100101101",36836 => "0000000100101101",
36837 => "0000000100101101",36838 => "0000000100101101",
36839 => "0000000100101101",36840 => "0000000000000011",
36841 => "0000000000000011",36842 => "0000000000000011",
36843 => "0000000000000011",36844 => "0000000000000011",
36845 => "0000000000000011",36846 => "0000000000000011",
36847 => "0000000000000011",36848 => "0000000000000011",
36849 => "0000000000000011",36850 => "0000000000000011",
36851 => "0000000000000011",36852 => "0000000000000011",
36853 => "0000000000000011",36854 => "0000000000000011",
36855 => "0000000000000011",36856 => "0000000000000011",
36857 => "0000000000000011",36858 => "0000000000000011",
36859 => "0000000000000011",36860 => "0000000000000011",
36861 => "0000000000000011",36862 => "0000000000000011",
36863 => "0000000000000011",36864 => "0000000010000111",
36865 => "0000000001111010",36866 => "0000000001101111",
36867 => "0000000000000001",36868 => "0000000001011011",
36869 => "0000000001010010",36870 => "0000000001001010",
36871 => "0000000001000011",36872 => "0000000000111101",
36873 => "0000000000110111",36874 => "0000000001111010",
36875 => "0000000001111001",36876 => "0000000000001100",
36877 => "0000000001110111",36878 => "0000000001110110",
36879 => "0000000001110100",36880 => "0000000001110011",
36881 => "0000000001110010",36882 => "0000000001110001",
36883 => "0000000001110000",36884 => "0000000001101111",
36885 => "0000000000001011",36886 => "0000000001101101",
36887 => "0000000001101100",36888 => "0000000001101010",
36889 => "0000000001101001",36890 => "0000000001101000",
36891 => "0000000001100111",36892 => "0000000001100110",
36893 => "0000000001100101",36894 => "0000000000000001",
36895 => "0000000001100011",36896 => "0000000001100010",
36897 => "0000000001100001",36898 => "0000000001100000",
36899 => "0000000001011111",36900 => "0000000001011110",
36901 => "0000000001011101",36902 => "0000000001011101",
36903 => "0000000001011100",36904 => "0000000001011011",
36905 => "0000000000001001",36906 => "0000000001011001",
36907 => "0000000001011000",36908 => "0000000001010111",
36909 => "0000000001010110",36910 => "0000000001010101",
36911 => "0000000001010101",36912 => "0000000001010100",
36913 => "0000000001010011",36914 => "0000000001010010",
36915 => "0000000001010001",36916 => "0000000000001000",
36917 => "0000000000001000",36918 => "0000000001001111",
36919 => "0000000001001110",36920 => "0000000001001101",
36921 => "0000000001001101",36922 => "0000000001001100",
36923 => "0000000001001011",36924 => "0000000001001010",
36925 => "0000000001001010",36926 => "0000000001001001",
36927 => "0000000001001000",36928 => "0000000001000111",
36929 => "0000000001000111",36930 => "0000000000000111",
36931 => "0000000001000101",36932 => "0000000001000101",
36933 => "0000000001000100",36934 => "0000000001000011",
36935 => "0000000001000011",36936 => "0000000001000010",
36937 => "0000000001000001",36938 => "0000000001000001",
36939 => "0000000001000000",36940 => "0000000000111111",
36941 => "0000000000111111",36942 => "0000000000111110",
36943 => "0000000000111101",36944 => "0000000000111101",
36945 => "0000000000000110",36946 => "0000000000000110",
36947 => "0000000000111011",36948 => "0000000000111010",
36949 => "0000000000111010",36950 => "0000000000111001",
36951 => "0000000000111001",36952 => "0000000000111000",
36953 => "0000000000111000",36954 => "0000000000110111",
36955 => "0000000000110110",36956 => "0000000000110110",
36957 => "0000000000110101",36958 => "0000000000110101",
36959 => "0000000000110100",36960 => "0000000000110100",
36961 => "0000000000110011",36962 => "0000000000110011",
36963 => "0000000000000101",36964 => "0000000001111010",
36965 => "0000000001111010",36966 => "0000000001111010",
36967 => "0000000001111010",36968 => "0000000001111010",
36969 => "0000000001111010",36970 => "0000000001111010",
36971 => "0000000001111010",36972 => "0000000001111001",
36973 => "0000000001111001",36974 => "0000000001111001",
36975 => "0000000001111001",36976 => "0000000001111001",
36977 => "0000000001111001",36978 => "0000000001111001",
36979 => "0000000001111001",36980 => "0000000001111001",
36981 => "0000000000001100",36982 => "0000000000001100",
36983 => "0000000000001100",36984 => "0000000000001100",
36985 => "0000000000001100",36986 => "0000000000001100",
36987 => "0000000000001100",36988 => "0000000000001100",
36989 => "0000000001110111",36990 => "0000000001110111",
36991 => "0000000001110111",36992 => "0000000001110111",
36993 => "0000000001110111",36994 => "0000000001110111",
36995 => "0000000001110111",36996 => "0000000001110111",
36997 => "0000000001110110",36998 => "0000000001110110",
36999 => "0000000001110110",37000 => "0000000001110110",
37001 => "0000000001110110",37002 => "0000000001110110",
37003 => "0000000001110110",37004 => "0000000001110110",
37005 => "0000000001110110",37006 => "0000000001110101",
37007 => "0000000001110101",37008 => "0000000001110101",
37009 => "0000000001110101",37010 => "0000000001110101",
37011 => "0000000001110101",37012 => "0000000001110101",
37013 => "0000000001110101",37014 => "0000000001110100",
37015 => "0000000001110100",37016 => "0000000001110100",
37017 => "0000000001110100",37018 => "0000000001110100",
37019 => "0000000001110100",37020 => "0000000001110100",
37021 => "0000000001110100",37022 => "0000000001110100",
37023 => "0000000001110011",37024 => "0000000001110011",
37025 => "0000000001110011",37026 => "0000000001110011",
37027 => "0000000001110011",37028 => "0000000001110011",
37029 => "0000000001110011",37030 => "0000000001110011",
37031 => "0000000001110011",37032 => "0000000001110010",
37033 => "0000000001110010",37034 => "0000000001110010",
37035 => "0000000001110010",37036 => "0000000001110010",
37037 => "0000000001110010",37038 => "0000000001110010",
37039 => "0000000001110010",37040 => "0000000001110001",
37041 => "0000000001110001",37042 => "0000000001110001",
37043 => "0000000001110001",37044 => "0000000001110001",
37045 => "0000000001110001",37046 => "0000000001110001",
37047 => "0000000001110001",37048 => "0000000001110001",
37049 => "0000000001110000",37050 => "0000000001110000",
37051 => "0000000001110000",37052 => "0000000001110000",
37053 => "0000000001110000",37054 => "0000000001110000",
37055 => "0000000001110000",37056 => "0000000001110000",
37057 => "0000000001110000",37058 => "0000000001101111",
37059 => "0000000001101111",37060 => "0000000001101111",
37061 => "0000000001101111",37062 => "0000000001101111",
37063 => "0000000001101111",37064 => "0000000001101111",
37065 => "0000000001101111",37066 => "0000000001101111",
37067 => "0000000000001011",37068 => "0000000000001011",
37069 => "0000000000001011",37070 => "0000000000001011",
37071 => "0000000000001011",37072 => "0000000000001011",
37073 => "0000000000001011",37074 => "0000000000001011",
37075 => "0000000000001011",37076 => "0000000001101101",
37077 => "0000000001101101",37078 => "0000000001101101",
37079 => "0000000001101101",37080 => "0000000001101101",
37081 => "0000000001101101",37082 => "0000000001101101",
37083 => "0000000001101101",37084 => "0000000001101101",
37085 => "0000000001101101",37086 => "0000000001101100",
37087 => "0000000001101100",37088 => "0000000001101100",
37089 => "0000000001101100",37090 => "0000000001101100",
37091 => "0000000001101100",37092 => "0000000001101100",
37093 => "0000000001101100",37094 => "0000000001101100",
37095 => "0000000001101011",37096 => "0000000001101011",
37097 => "0000000001101011",37098 => "0000000001101011",
37099 => "0000000001101011",37100 => "0000000001101011",
37101 => "0000000001101011",37102 => "0000000001101011",
37103 => "0000000001101011",37104 => "0000000001101010",
37105 => "0000000001101010",37106 => "0000000001101010",
37107 => "0000000001101010",37108 => "0000000001101010",
37109 => "0000000001101010",37110 => "0000000001101010",
37111 => "0000000001101010",37112 => "0000000001101010",
37113 => "0000000001101010",37114 => "0000000001101001",
37115 => "0000000001101001",37116 => "0000000001101001",
37117 => "0000000001101001",37118 => "0000000001101001",
37119 => "0000000001101001",37120 => "0000000001101001",
37121 => "0000000001101001",37122 => "0000000001101001",
37123 => "0000000001101000",37124 => "0000000001101000",
37125 => "0000000001101000",37126 => "0000000001101000",
37127 => "0000000001101000",37128 => "0000000001101000",
37129 => "0000000001101000",37130 => "0000000001101000",
37131 => "0000000001101000",37132 => "0000000001101000",
37133 => "0000000001100111",37134 => "0000000001100111",
37135 => "0000000001100111",37136 => "0000000001100111",
37137 => "0000000001100111",37138 => "0000000001100111",
37139 => "0000000001100111",37140 => "0000000001100111",
37141 => "0000000001100111",37142 => "0000000001100110",
37143 => "0000000001100110",37144 => "0000000001100110",
37145 => "0000000001100110",37146 => "0000000001100110",
37147 => "0000000001100110",37148 => "0000000001100110",
37149 => "0000000001100110",37150 => "0000000001100110",
37151 => "0000000001100110",37152 => "0000000001100101",
37153 => "0000000001100101",37154 => "0000000001100101",
37155 => "0000000001100101",37156 => "0000000001100101",
37157 => "0000000001100101",37158 => "0000000001100101",
37159 => "0000000001100101",37160 => "0000000001100101",
37161 => "0000000001100101",37162 => "0000000000000001",
37163 => "0000000000000001",37164 => "0000000000000001",
37165 => "0000000000000001",37166 => "0000000000000001",
37167 => "0000000000000001",37168 => "0000000000000001",
37169 => "0000000000000001",37170 => "0000000000000001",
37171 => "0000000000000001",37172 => "0000000001100011",
37173 => "0000000001100011",37174 => "0000000001100011",
37175 => "0000000001100011",37176 => "0000000001100011",
37177 => "0000000001100011",37178 => "0000000001100011",
37179 => "0000000001100011",37180 => "0000000001100011",
37181 => "0000000001100011",37182 => "0000000001100010",
37183 => "0000000001100010",37184 => "0000000001100010",
37185 => "0000000001100010",37186 => "0000000001100010",
37187 => "0000000001100010",37188 => "0000000001100010",
37189 => "0000000001100010",37190 => "0000000001100010",
37191 => "0000000001100010",37192 => "0000000001100001",
37193 => "0000000001100001",37194 => "0000000001100001",
37195 => "0000000001100001",37196 => "0000000001100001",
37197 => "0000000001100001",37198 => "0000000001100001",
37199 => "0000000001100001",37200 => "0000000001100001",
37201 => "0000000001100001",37202 => "0000000001100001",
37203 => "0000000001100000",37204 => "0000000001100000",
37205 => "0000000001100000",37206 => "0000000001100000",
37207 => "0000000001100000",37208 => "0000000001100000",
37209 => "0000000001100000",37210 => "0000000001100000",
37211 => "0000000001100000",37212 => "0000000001100000",
37213 => "0000000001011111",37214 => "0000000001011111",
37215 => "0000000001011111",37216 => "0000000001011111",
37217 => "0000000001011111",37218 => "0000000001011111",
37219 => "0000000001011111",37220 => "0000000001011111",
37221 => "0000000001011111",37222 => "0000000001011111",
37223 => "0000000001011111",37224 => "0000000001011110",
37225 => "0000000001011110",37226 => "0000000001011110",
37227 => "0000000001011110",37228 => "0000000001011110",
37229 => "0000000001011110",37230 => "0000000001011110",
37231 => "0000000001011110",37232 => "0000000001011110",
37233 => "0000000001011110",37234 => "0000000001011101",
37235 => "0000000001011101",37236 => "0000000001011101",
37237 => "0000000001011101",37238 => "0000000001011101",
37239 => "0000000001011101",37240 => "0000000001011101",
37241 => "0000000001011101",37242 => "0000000001011101",
37243 => "0000000001011101",37244 => "0000000001011101",
37245 => "0000000001011100",37246 => "0000000001011100",
37247 => "0000000001011100",37248 => "0000000001011100",
37249 => "0000000001011100",37250 => "0000000001011100",
37251 => "0000000001011100",37252 => "0000000001011100",
37253 => "0000000001011100",37254 => "0000000001011100",
37255 => "0000000001011100",37256 => "0000000001011011",
37257 => "0000000001011011",37258 => "0000000001011011",
37259 => "0000000001011011",37260 => "0000000001011011",
37261 => "0000000001011011",37262 => "0000000001011011",
37263 => "0000000001011011",37264 => "0000000001011011",
37265 => "0000000001011011",37266 => "0000000001011011",
37267 => "0000000000001001",37268 => "0000000000001001",
37269 => "0000000000001001",37270 => "0000000000001001",
37271 => "0000000000001001",37272 => "0000000000001001",
37273 => "0000000000001001",37274 => "0000000000001001",
37275 => "0000000000001001",37276 => "0000000000001001",
37277 => "0000000000001001",37278 => "0000000001011001",
37279 => "0000000001011001",37280 => "0000000001011001",
37281 => "0000000001011001",37282 => "0000000001011001",
37283 => "0000000001011001",37284 => "0000000001011001",
37285 => "0000000001011001",37286 => "0000000001011001",
37287 => "0000000001011001",37288 => "0000000001011001",
37289 => "0000000001011000",37290 => "0000000001011000",
37291 => "0000000001011000",37292 => "0000000001011000",
37293 => "0000000001011000",37294 => "0000000001011000",
37295 => "0000000001011000",37296 => "0000000001011000",
37297 => "0000000001011000",37298 => "0000000001011000",
37299 => "0000000001011000",37300 => "0000000001011000",
37301 => "0000000001010111",37302 => "0000000001010111",
37303 => "0000000001010111",37304 => "0000000001010111",
37305 => "0000000001010111",37306 => "0000000001010111",
37307 => "0000000001010111",37308 => "0000000001010111",
37309 => "0000000001010111",37310 => "0000000001010111",
37311 => "0000000001010111",37312 => "0000000001010110",
37313 => "0000000001010110",37314 => "0000000001010110",
37315 => "0000000001010110",37316 => "0000000001010110",
37317 => "0000000001010110",37318 => "0000000001010110",
37319 => "0000000001010110",37320 => "0000000001010110",
37321 => "0000000001010110",37322 => "0000000001010110",
37323 => "0000000001010110",37324 => "0000000001010101",
37325 => "0000000001010101",37326 => "0000000001010101",
37327 => "0000000001010101",37328 => "0000000001010101",
37329 => "0000000001010101",37330 => "0000000001010101",
37331 => "0000000001010101",37332 => "0000000001010101",
37333 => "0000000001010101",37334 => "0000000001010101",
37335 => "0000000001010101",37336 => "0000000001010100",
37337 => "0000000001010100",37338 => "0000000001010100",
37339 => "0000000001010100",37340 => "0000000001010100",
37341 => "0000000001010100",37342 => "0000000001010100",
37343 => "0000000001010100",37344 => "0000000001010100",
37345 => "0000000001010100",37346 => "0000000001010100",
37347 => "0000000001010011",37348 => "0000000001010011",
37349 => "0000000001010011",37350 => "0000000001010011",
37351 => "0000000001010011",37352 => "0000000001010011",
37353 => "0000000001010011",37354 => "0000000001010011",
37355 => "0000000001010011",37356 => "0000000001010011",
37357 => "0000000001010011",37358 => "0000000001010011",
37359 => "0000000001010010",37360 => "0000000001010010",
37361 => "0000000001010010",37362 => "0000000001010010",
37363 => "0000000001010010",37364 => "0000000001010010",
37365 => "0000000001010010",37366 => "0000000001010010",
37367 => "0000000001010010",37368 => "0000000001010010",
37369 => "0000000001010010",37370 => "0000000001010010",
37371 => "0000000001010010",37372 => "0000000001010001",
37373 => "0000000001010001",37374 => "0000000001010001",
37375 => "0000000001010001",37376 => "0000000001010001",
37377 => "0000000001010001",37378 => "0000000001010001",
37379 => "0000000001010001",37380 => "0000000001010001",
37381 => "0000000001010001",37382 => "0000000001010001",
37383 => "0000000001010001",37384 => "0000000000001000",
37385 => "0000000000001000",37386 => "0000000000001000",
37387 => "0000000000001000",37388 => "0000000000001000",
37389 => "0000000000001000",37390 => "0000000000001000",
37391 => "0000000000001000",37392 => "0000000000001000",
37393 => "0000000000001000",37394 => "0000000000001000",
37395 => "0000000000001000",37396 => "0000000001001111",
37397 => "0000000001001111",37398 => "0000000001001111",
37399 => "0000000001001111",37400 => "0000000001001111",
37401 => "0000000001001111",37402 => "0000000001001111",
37403 => "0000000001001111",37404 => "0000000001001111",
37405 => "0000000001001111",37406 => "0000000001001111",
37407 => "0000000001001111",37408 => "0000000001001111",
37409 => "0000000001001110",37410 => "0000000001001110",
37411 => "0000000001001110",37412 => "0000000001001110",
37413 => "0000000001001110",37414 => "0000000001001110",
37415 => "0000000001001110",37416 => "0000000001001110",
37417 => "0000000001001110",37418 => "0000000001001110",
37419 => "0000000001001110",37420 => "0000000001001110",
37421 => "0000000001001110",37422 => "0000000001001101",
37423 => "0000000001001101",37424 => "0000000001001101",
37425 => "0000000001001101",37426 => "0000000001001101",
37427 => "0000000001001101",37428 => "0000000001001101",
37429 => "0000000001001101",37430 => "0000000001001101",
37431 => "0000000001001101",37432 => "0000000001001101",
37433 => "0000000001001101",37434 => "0000000001001101",
37435 => "0000000001001100",37436 => "0000000001001100",
37437 => "0000000001001100",37438 => "0000000001001100",
37439 => "0000000001001100",37440 => "0000000001001100",
37441 => "0000000001001100",37442 => "0000000001001100",
37443 => "0000000001001100",37444 => "0000000001001100",
37445 => "0000000001001100",37446 => "0000000001001100",
37447 => "0000000001001100",37448 => "0000000001001011",
37449 => "0000000001001011",37450 => "0000000001001011",
37451 => "0000000001001011",37452 => "0000000001001011",
37453 => "0000000001001011",37454 => "0000000001001011",
37455 => "0000000001001011",37456 => "0000000001001011",
37457 => "0000000001001011",37458 => "0000000001001011",
37459 => "0000000001001011",37460 => "0000000001001011",
37461 => "0000000001001010",37462 => "0000000001001010",
37463 => "0000000001001010",37464 => "0000000001001010",
37465 => "0000000001001010",37466 => "0000000001001010",
37467 => "0000000001001010",37468 => "0000000001001010",
37469 => "0000000001001010",37470 => "0000000001001010",
37471 => "0000000001001010",37472 => "0000000001001010",
37473 => "0000000001001010",37474 => "0000000001001010",
37475 => "0000000001001001",37476 => "0000000001001001",
37477 => "0000000001001001",37478 => "0000000001001001",
37479 => "0000000001001001",37480 => "0000000001001001",
37481 => "0000000001001001",37482 => "0000000001001001",
37483 => "0000000001001001",37484 => "0000000001001001",
37485 => "0000000001001001",37486 => "0000000001001001",
37487 => "0000000001001001",37488 => "0000000001001001",
37489 => "0000000001001000",37490 => "0000000001001000",
37491 => "0000000001001000",37492 => "0000000001001000",
37493 => "0000000001001000",37494 => "0000000001001000",
37495 => "0000000001001000",37496 => "0000000001001000",
37497 => "0000000001001000",37498 => "0000000001001000",
37499 => "0000000001001000",37500 => "0000000001001000",
37501 => "0000000001001000",37502 => "0000000001001000",
37503 => "0000000001000111",37504 => "0000000001000111",
37505 => "0000000001000111",37506 => "0000000001000111",
37507 => "0000000001000111",37508 => "0000000001000111",
37509 => "0000000001000111",37510 => "0000000001000111",
37511 => "0000000001000111",37512 => "0000000001000111",
37513 => "0000000001000111",37514 => "0000000001000111",
37515 => "0000000001000111",37516 => "0000000001000111",
37517 => "0000000000000111",37518 => "0000000000000111",
37519 => "0000000000000111",37520 => "0000000000000111",
37521 => "0000000000000111",37522 => "0000000000000111",
37523 => "0000000000000111",37524 => "0000000000000111",
37525 => "0000000000000111",37526 => "0000000000000111",
37527 => "0000000000000111",37528 => "0000000000000111",
37529 => "0000000000000111",37530 => "0000000000000111",
37531 => "0000000001000101",37532 => "0000000001000101",
37533 => "0000000001000101",37534 => "0000000001000101",
37535 => "0000000001000101",37536 => "0000000001000101",
37537 => "0000000001000101",37538 => "0000000001000101",
37539 => "0000000001000101",37540 => "0000000001000101",
37541 => "0000000001000101",37542 => "0000000001000101",
37543 => "0000000001000101",37544 => "0000000001000101",
37545 => "0000000001000100",37546 => "0000000001000100",
37547 => "0000000001000100",37548 => "0000000001000100",
37549 => "0000000001000100",37550 => "0000000001000100",
37551 => "0000000001000100",37552 => "0000000001000100",
37553 => "0000000001000100",37554 => "0000000001000100",
37555 => "0000000001000100",37556 => "0000000001000100",
37557 => "0000000001000100",37558 => "0000000001000100",
37559 => "0000000001000100",37560 => "0000000001000011",
37561 => "0000000001000011",37562 => "0000000001000011",
37563 => "0000000001000011",37564 => "0000000001000011",
37565 => "0000000001000011",37566 => "0000000001000011",
37567 => "0000000001000011",37568 => "0000000001000011",
37569 => "0000000001000011",37570 => "0000000001000011",
37571 => "0000000001000011",37572 => "0000000001000011",
37573 => "0000000001000011",37574 => "0000000001000011",
37575 => "0000000001000010",37576 => "0000000001000010",
37577 => "0000000001000010",37578 => "0000000001000010",
37579 => "0000000001000010",37580 => "0000000001000010",
37581 => "0000000001000010",37582 => "0000000001000010",
37583 => "0000000001000010",37584 => "0000000001000010",
37585 => "0000000001000010",37586 => "0000000001000010",
37587 => "0000000001000010",37588 => "0000000001000010",
37589 => "0000000001000010",37590 => "0000000001000001",
37591 => "0000000001000001",37592 => "0000000001000001",
37593 => "0000000001000001",37594 => "0000000001000001",
37595 => "0000000001000001",37596 => "0000000001000001",
37597 => "0000000001000001",37598 => "0000000001000001",
37599 => "0000000001000001",37600 => "0000000001000001",
37601 => "0000000001000001",37602 => "0000000001000001",
37603 => "0000000001000001",37604 => "0000000001000001",
37605 => "0000000001000001",37606 => "0000000001000000",
37607 => "0000000001000000",37608 => "0000000001000000",
37609 => "0000000001000000",37610 => "0000000001000000",
37611 => "0000000001000000",37612 => "0000000001000000",
37613 => "0000000001000000",37614 => "0000000001000000",
37615 => "0000000001000000",37616 => "0000000001000000",
37617 => "0000000001000000",37618 => "0000000001000000",
37619 => "0000000001000000",37620 => "0000000001000000",
37621 => "0000000000111111",37622 => "0000000000111111",
37623 => "0000000000111111",37624 => "0000000000111111",
37625 => "0000000000111111",37626 => "0000000000111111",
37627 => "0000000000111111",37628 => "0000000000111111",
37629 => "0000000000111111",37630 => "0000000000111111",
37631 => "0000000000111111",37632 => "0000000000111111",
37633 => "0000000000111111",37634 => "0000000000111111",
37635 => "0000000000111111",37636 => "0000000000111111",
37637 => "0000000000111110",37638 => "0000000000111110",
37639 => "0000000000111110",37640 => "0000000000111110",
37641 => "0000000000111110",37642 => "0000000000111110",
37643 => "0000000000111110",37644 => "0000000000111110",
37645 => "0000000000111110",37646 => "0000000000111110",
37647 => "0000000000111110",37648 => "0000000000111110",
37649 => "0000000000111110",37650 => "0000000000111110",
37651 => "0000000000111110",37652 => "0000000000111110",
37653 => "0000000000111101",37654 => "0000000000111101",
37655 => "0000000000111101",37656 => "0000000000111101",
37657 => "0000000000111101",37658 => "0000000000111101",
37659 => "0000000000111101",37660 => "0000000000111101",
37661 => "0000000000111101",37662 => "0000000000111101",
37663 => "0000000000111101",37664 => "0000000000111101",
37665 => "0000000000111101",37666 => "0000000000111101",
37667 => "0000000000111101",37668 => "0000000000111101",
37669 => "0000000000111101",37670 => "0000000000000110",
37671 => "0000000000000110",37672 => "0000000000000110",
37673 => "0000000000000110",37674 => "0000000000000110",
37675 => "0000000000000110",37676 => "0000000000000110",
37677 => "0000000000000110",37678 => "0000000000000110",
37679 => "0000000000000110",37680 => "0000000000000110",
37681 => "0000000000000110",37682 => "0000000000000110",
37683 => "0000000000000110",37684 => "0000000000000110",
37685 => "0000000000000110",37686 => "0000000000111011",
37687 => "0000000000111011",37688 => "0000000000111011",
37689 => "0000000000111011",37690 => "0000000000111011",
37691 => "0000000000111011",37692 => "0000000000111011",
37693 => "0000000000111011",37694 => "0000000000111011",
37695 => "0000000000111011",37696 => "0000000000111011",
37697 => "0000000000111011",37698 => "0000000000111011",
37699 => "0000000000111011",37700 => "0000000000111011",
37701 => "0000000000111011",37702 => "0000000000111011",
37703 => "0000000000111010",37704 => "0000000000111010",
37705 => "0000000000111010",37706 => "0000000000111010",
37707 => "0000000000111010",37708 => "0000000000111010",
37709 => "0000000000111010",37710 => "0000000000111010",
37711 => "0000000000111010",37712 => "0000000000111010",
37713 => "0000000000111010",37714 => "0000000000111010",
37715 => "0000000000111010",37716 => "0000000000111010",
37717 => "0000000000111010",37718 => "0000000000111010",
37719 => "0000000000111010",37720 => "0000000000111001",
37721 => "0000000000111001",37722 => "0000000000111001",
37723 => "0000000000111001",37724 => "0000000000111001",
37725 => "0000000000111001",37726 => "0000000000111001",
37727 => "0000000000111001",37728 => "0000000000111001",
37729 => "0000000000111001",37730 => "0000000000111001",
37731 => "0000000000111001",37732 => "0000000000111001",
37733 => "0000000000111001",37734 => "0000000000111001",
37735 => "0000000000111001",37736 => "0000000000111001",
37737 => "0000000000111001",37738 => "0000000000111000",
37739 => "0000000000111000",37740 => "0000000000111000",
37741 => "0000000000111000",37742 => "0000000000111000",
37743 => "0000000000111000",37744 => "0000000000111000",
37745 => "0000000000111000",37746 => "0000000000111000",
37747 => "0000000000111000",37748 => "0000000000111000",
37749 => "0000000000111000",37750 => "0000000000111000",
37751 => "0000000000111000",37752 => "0000000000111000",
37753 => "0000000000111000",37754 => "0000000000111000",
37755 => "0000000000111000",37756 => "0000000000110111",
37757 => "0000000000110111",37758 => "0000000000110111",
37759 => "0000000000110111",37760 => "0000000000110111",
37761 => "0000000000110111",37762 => "0000000000110111",
37763 => "0000000000110111",37764 => "0000000000110111",
37765 => "0000000000110111",37766 => "0000000000110111",
37767 => "0000000000110111",37768 => "0000000000110111",
37769 => "0000000000110111",37770 => "0000000000110111",
37771 => "0000000000110111",37772 => "0000000000110111",
37773 => "0000000000110111",37774 => "0000000000110110",
37775 => "0000000000110110",37776 => "0000000000110110",
37777 => "0000000000110110",37778 => "0000000000110110",
37779 => "0000000000110110",37780 => "0000000000110110",
37781 => "0000000000110110",37782 => "0000000000110110",
37783 => "0000000000110110",37784 => "0000000000110110",
37785 => "0000000000110110",37786 => "0000000000110110",
37787 => "0000000000110110",37788 => "0000000000110110",
37789 => "0000000000110110",37790 => "0000000000110110",
37791 => "0000000000110110",37792 => "0000000000110110",
37793 => "0000000000110101",37794 => "0000000000110101",
37795 => "0000000000110101",37796 => "0000000000110101",
37797 => "0000000000110101",37798 => "0000000000110101",
37799 => "0000000000110101",37800 => "0000000000110101",
37801 => "0000000000110101",37802 => "0000000000110101",
37803 => "0000000000110101",37804 => "0000000000110101",
37805 => "0000000000110101",37806 => "0000000000110101",
37807 => "0000000000110101",37808 => "0000000000110101",
37809 => "0000000000110101",37810 => "0000000000110101",
37811 => "0000000000110100",37812 => "0000000000110100",
37813 => "0000000000110100",37814 => "0000000000110100",
37815 => "0000000000110100",37816 => "0000000000110100",
37817 => "0000000000110100",37818 => "0000000000110100",
37819 => "0000000000110100",37820 => "0000000000110100",
37821 => "0000000000110100",37822 => "0000000000110100",
37823 => "0000000000110100",37824 => "0000000000110100",
37825 => "0000000000110100",37826 => "0000000000110100",
37827 => "0000000000110100",37828 => "0000000000110100",
37829 => "0000000000110100",37830 => "0000000000110100",
37831 => "0000000000110011",37832 => "0000000000110011",
37833 => "0000000000110011",37834 => "0000000000110011",
37835 => "0000000000110011",37836 => "0000000000110011",
37837 => "0000000000110011",37838 => "0000000000110011",
37839 => "0000000000110011",37840 => "0000000000110011",
37841 => "0000000000110011",37842 => "0000000000110011",
37843 => "0000000000110011",37844 => "0000000000110011",
37845 => "0000000000110011",37846 => "0000000000110011",
37847 => "0000000000110011",37848 => "0000000000110011",
37849 => "0000000000110011",37850 => "0000000000000101",
37851 => "0000000000000101",37852 => "0000000000000101",
37853 => "0000000000000101",37854 => "0000000000000101",
37855 => "0000000000000101",37856 => "0000000000000101",
37857 => "0000000000000101",37858 => "0000000000000101",
37859 => "0000000000000101",37860 => "0000000000000101",
37861 => "0000000000000101",37862 => "0000000000000101",
37863 => "0000000000000101",37864 => "0000000001111010",
37865 => "0000000001111010",37866 => "0000000001111010",
37867 => "0000000001111010",37868 => "0000000001111010",
37869 => "0000000001111010",37870 => "0000000001111010",
37871 => "0000000001111010",37872 => "0000000001111010",
37873 => "0000000001111010",37874 => "0000000001111010",
37875 => "0000000001111010",37876 => "0000000001111010",
37877 => "0000000001111010",37878 => "0000000001111010",
37879 => "0000000001111010",37880 => "0000000001111010",
37881 => "0000000001111010",37882 => "0000000001111010",
37883 => "0000000001111010",37884 => "0000000001111010",
37885 => "0000000001111010",37886 => "0000000001111010",
37887 => "0000000001111010",37888 => "0000000001111010",
37889 => "0000000001111010",37890 => "0000000001111010",
37891 => "0000000001111010",37892 => "0000000001111010",
37893 => "0000000001111010",37894 => "0000000001111010",
37895 => "0000000001111010",37896 => "0000000001111010",
37897 => "0000000001111010",37898 => "0000000001111010",
37899 => "0000000001111010",37900 => "0000000001111010",
37901 => "0000000001111010",37902 => "0000000001111010",
37903 => "0000000001111010",37904 => "0000000001111010",
37905 => "0000000001111010",37906 => "0000000001111010",
37907 => "0000000001111010",37908 => "0000000001111010",
37909 => "0000000001111010",37910 => "0000000001111010",
37911 => "0000000001111010",37912 => "0000000001111010",
37913 => "0000000001111010",37914 => "0000000001111010",
37915 => "0000000001111010",37916 => "0000000001111010",
37917 => "0000000001111010",37918 => "0000000001111010",
37919 => "0000000001111010",37920 => "0000000001111010",
37921 => "0000000001111010",37922 => "0000000001111010",
37923 => "0000000001111010",37924 => "0000000001111010",
37925 => "0000000001111010",37926 => "0000000001111010",
37927 => "0000000001111010",37928 => "0000000001111010",
37929 => "0000000001111010",37930 => "0000000001111010",
37931 => "0000000001111010",37932 => "0000000001111010",
37933 => "0000000001111010",37934 => "0000000001111010",
37935 => "0000000001111010",37936 => "0000000001111010",
37937 => "0000000001111010",37938 => "0000000001111010",
37939 => "0000000001111010",37940 => "0000000001111010",
37941 => "0000000001111010",37942 => "0000000001111010",
37943 => "0000000001111001",37944 => "0000000001111001",
37945 => "0000000001111001",37946 => "0000000001111001",
37947 => "0000000001111001",37948 => "0000000001111001",
37949 => "0000000001111001",37950 => "0000000001111001",
37951 => "0000000001111001",37952 => "0000000001111001",
37953 => "0000000001111001",37954 => "0000000001111001",
37955 => "0000000001111001",37956 => "0000000001111001",
37957 => "0000000001111001",37958 => "0000000001111001",
37959 => "0000000001111001",37960 => "0000000001111001",
37961 => "0000000001111001",37962 => "0000000001111001",
37963 => "0000000001111001",37964 => "0000000001111001",
37965 => "0000000001111001",37966 => "0000000001111001",
37967 => "0000000001111001",37968 => "0000000001111001",
37969 => "0000000001111001",37970 => "0000000001111001",
37971 => "0000000001111001",37972 => "0000000001111001",
37973 => "0000000001111001",37974 => "0000000001111001",
37975 => "0000000001111001",37976 => "0000000001111001",
37977 => "0000000001111001",37978 => "0000000001111001",
37979 => "0000000001111001",37980 => "0000000001111001",
37981 => "0000000001111001",37982 => "0000000001111001",
37983 => "0000000001111001",37984 => "0000000001111001",
37985 => "0000000001111001",37986 => "0000000001111001",
37987 => "0000000001111001",37988 => "0000000001111001",
37989 => "0000000001111001",37990 => "0000000001111001",
37991 => "0000000001111001",37992 => "0000000001111001",
37993 => "0000000001111001",37994 => "0000000001111001",
37995 => "0000000001111001",37996 => "0000000001111001",
37997 => "0000000001111001",37998 => "0000000001111001",
37999 => "0000000001111001",38000 => "0000000001111001",
38001 => "0000000001111001",38002 => "0000000001111001",
38003 => "0000000001111001",38004 => "0000000001111001",
38005 => "0000000001111001",38006 => "0000000001111001",
38007 => "0000000001111001",38008 => "0000000001111001",
38009 => "0000000001111001",38010 => "0000000001111001",
38011 => "0000000001111001",38012 => "0000000001111001",
38013 => "0000000001111001",38014 => "0000000001111001",
38015 => "0000000001111001",38016 => "0000000001111001",
38017 => "0000000001111001",38018 => "0000000001111001",
38019 => "0000000001111001",38020 => "0000000001111001",
38021 => "0000000001111001",38022 => "0000000001111001",
38023 => "0000000001111001",38024 => "0000000001111001",
38025 => "0000000001111001",38026 => "0000000000001100",
38027 => "0000000000001100",38028 => "0000000000001100",
38029 => "0000000000001100",38030 => "0000000000001100",
38031 => "0000000000001100",38032 => "0000000000001100",
38033 => "0000000000001100",38034 => "0000000000001100",
38035 => "0000000000001100",38036 => "0000000000001100",
38037 => "0000000000001100",38038 => "0000000000001100",
38039 => "0000000000001100",38040 => "0000000000001100",
38041 => "0000000000001100",38042 => "0000000000001100",
38043 => "0000000000001100",38044 => "0000000000001100",
38045 => "0000000000001100",38046 => "0000000000001100",
38047 => "0000000000001100",38048 => "0000000000001100",
38049 => "0000000000001100",38050 => "0000000000001100",
38051 => "0000000000001100",38052 => "0000000000001100",
38053 => "0000000000001100",38054 => "0000000000001100",
38055 => "0000000000001100",38056 => "0000000000001100",
38057 => "0000000000001100",38058 => "0000000000001100",
38059 => "0000000000001100",38060 => "0000000000001100",
38061 => "0000000000001100",38062 => "0000000000001100",
38063 => "0000000000001100",38064 => "0000000000001100",
38065 => "0000000000001100",38066 => "0000000000001100",
38067 => "0000000000001100",38068 => "0000000000001100",
38069 => "0000000000001100",38070 => "0000000000001100",
38071 => "0000000000001100",38072 => "0000000000001100",
38073 => "0000000000001100",38074 => "0000000000001100",
38075 => "0000000000001100",38076 => "0000000000001100",
38077 => "0000000000001100",38078 => "0000000000001100",
38079 => "0000000000001100",38080 => "0000000000001100",
38081 => "0000000000001100",38082 => "0000000000001100",
38083 => "0000000000001100",38084 => "0000000000001100",
38085 => "0000000000001100",38086 => "0000000000001100",
38087 => "0000000000001100",38088 => "0000000000001100",
38089 => "0000000000001100",38090 => "0000000000001100",
38091 => "0000000000001100",38092 => "0000000000001100",
38093 => "0000000000001100",38094 => "0000000000001100",
38095 => "0000000000001100",38096 => "0000000000001100",
38097 => "0000000000001100",38098 => "0000000000001100",
38099 => "0000000000001100",38100 => "0000000000001100",
38101 => "0000000000001100",38102 => "0000000000001100",
38103 => "0000000000001100",38104 => "0000000000001100",
38105 => "0000000000001100",38106 => "0000000000001100",
38107 => "0000000000001100",38108 => "0000000000001100",
38109 => "0000000001110111",38110 => "0000000001110111",
38111 => "0000000001110111",38112 => "0000000001110111",
38113 => "0000000001110111",38114 => "0000000001110111",
38115 => "0000000001110111",38116 => "0000000001110111",
38117 => "0000000001110111",38118 => "0000000001110111",
38119 => "0000000001110111",38120 => "0000000001110111",
38121 => "0000000001110111",38122 => "0000000001110111",
38123 => "0000000001110111",38124 => "0000000001110111",
38125 => "0000000001110111",38126 => "0000000001110111",
38127 => "0000000001110111",38128 => "0000000001110111",
38129 => "0000000001110111",38130 => "0000000001110111",
38131 => "0000000001110111",38132 => "0000000001110111",
38133 => "0000000001110111",38134 => "0000000001110111",
38135 => "0000000001110111",38136 => "0000000001110111",
38137 => "0000000001110111",38138 => "0000000001110111",
38139 => "0000000001110111",38140 => "0000000001110111",
38141 => "0000000001110111",38142 => "0000000001110111",
38143 => "0000000001110111",38144 => "0000000001110111",
38145 => "0000000001110111",38146 => "0000000001110111",
38147 => "0000000001110111",38148 => "0000000001110111",
38149 => "0000000001110111",38150 => "0000000001110111",
38151 => "0000000001110111",38152 => "0000000001110111",
38153 => "0000000001110111",38154 => "0000000001110111",
38155 => "0000000001110111",38156 => "0000000001110111",
38157 => "0000000001110111",38158 => "0000000001110111",
38159 => "0000000001110111",38160 => "0000000001110111",
38161 => "0000000001110111",38162 => "0000000001110111",
38163 => "0000000001110111",38164 => "0000000001110111",
38165 => "0000000001110111",38166 => "0000000001110111",
38167 => "0000000001110111",38168 => "0000000001110111",
38169 => "0000000001110111",38170 => "0000000001110111",
38171 => "0000000001110111",38172 => "0000000001110111",
38173 => "0000000001110111",38174 => "0000000001110111",
38175 => "0000000001110111",38176 => "0000000001110111",
38177 => "0000000001110111",38178 => "0000000001110111",
38179 => "0000000001110111",38180 => "0000000001110111",
38181 => "0000000001110111",38182 => "0000000001110111",
38183 => "0000000001110111",38184 => "0000000001110111",
38185 => "0000000001110111",38186 => "0000000001110111",
38187 => "0000000001110111",38188 => "0000000001110111",
38189 => "0000000001110111",38190 => "0000000001110111",
38191 => "0000000001110111",38192 => "0000000001110111",
38193 => "0000000001110110",38194 => "0000000001110110",
38195 => "0000000001110110",38196 => "0000000001110110",
38197 => "0000000001110110",38198 => "0000000001110110",
38199 => "0000000001110110",38200 => "0000000001110110",
38201 => "0000000001110110",38202 => "0000000001110110",
38203 => "0000000001110110",38204 => "0000000001110110",
38205 => "0000000001110110",38206 => "0000000001110110",
38207 => "0000000001110110",38208 => "0000000001110110",
38209 => "0000000001110110",38210 => "0000000001110110",
38211 => "0000000001110110",38212 => "0000000001110110",
38213 => "0000000001110110",38214 => "0000000001110110",
38215 => "0000000001110110",38216 => "0000000001110110",
38217 => "0000000001110110",38218 => "0000000001110110",
38219 => "0000000001110110",38220 => "0000000001110110",
38221 => "0000000001110110",38222 => "0000000001110110",
38223 => "0000000001110110",38224 => "0000000001110110",
38225 => "0000000001110110",38226 => "0000000001110110",
38227 => "0000000001110110",38228 => "0000000001110110",
38229 => "0000000001110110",38230 => "0000000001110110",
38231 => "0000000001110110",38232 => "0000000001110110",
38233 => "0000000001110110",38234 => "0000000001110110",
38235 => "0000000001110110",38236 => "0000000001110110",
38237 => "0000000001110110",38238 => "0000000001110110",
38239 => "0000000001110110",38240 => "0000000001110110",
38241 => "0000000001110110",38242 => "0000000001110110",
38243 => "0000000001110110",38244 => "0000000001110110",
38245 => "0000000001110110",38246 => "0000000001110110",
38247 => "0000000001110110",38248 => "0000000001110110",
38249 => "0000000001110110",38250 => "0000000001110110",
38251 => "0000000001110110",38252 => "0000000001110110",
38253 => "0000000001110110",38254 => "0000000001110110",
38255 => "0000000001110110",38256 => "0000000001110110",
38257 => "0000000001110110",38258 => "0000000001110110",
38259 => "0000000001110110",38260 => "0000000001110110",
38261 => "0000000001110110",38262 => "0000000001110110",
38263 => "0000000001110110",38264 => "0000000001110110",
38265 => "0000000001110110",38266 => "0000000001110110",
38267 => "0000000001110110",38268 => "0000000001110110",
38269 => "0000000001110110",38270 => "0000000001110110",
38271 => "0000000001110110",38272 => "0000000001110110",
38273 => "0000000001110110",38274 => "0000000001110110",
38275 => "0000000001110110",38276 => "0000000001110110",
38277 => "0000000001110110",38278 => "0000000001110101",
38279 => "0000000001110101",38280 => "0000000001110101",
38281 => "0000000001110101",38282 => "0000000001110101",
38283 => "0000000001110101",38284 => "0000000001110101",
38285 => "0000000001110101",38286 => "0000000001110101",
38287 => "0000000001110101",38288 => "0000000001110101",
38289 => "0000000001110101",38290 => "0000000001110101",
38291 => "0000000001110101",38292 => "0000000001110101",
38293 => "0000000001110101",38294 => "0000000001110101",
38295 => "0000000001110101",38296 => "0000000001110101",
38297 => "0000000001110101",38298 => "0000000001110101",
38299 => "0000000001110101",38300 => "0000000001110101",
38301 => "0000000001110101",38302 => "0000000001110101",
38303 => "0000000001110101",38304 => "0000000001110101",
38305 => "0000000001110101",38306 => "0000000001110101",
38307 => "0000000001110101",38308 => "0000000001110101",
38309 => "0000000001110101",38310 => "0000000001110101",
38311 => "0000000001110101",38312 => "0000000001110101",
38313 => "0000000001110101",38314 => "0000000001110101",
38315 => "0000000001110101",38316 => "0000000001110101",
38317 => "0000000001110101",38318 => "0000000001110101",
38319 => "0000000001110101",38320 => "0000000001110101",
38321 => "0000000001110101",38322 => "0000000001110101",
38323 => "0000000001110101",38324 => "0000000001110101",
38325 => "0000000001110101",38326 => "0000000001110101",
38327 => "0000000001110101",38328 => "0000000001110101",
38329 => "0000000001110101",38330 => "0000000001110101",
38331 => "0000000001110101",38332 => "0000000001110101",
38333 => "0000000001110101",38334 => "0000000001110101",
38335 => "0000000001110101",38336 => "0000000001110101",
38337 => "0000000001110101",38338 => "0000000001110101",
38339 => "0000000001110101",38340 => "0000000001110101",
38341 => "0000000001110101",38342 => "0000000001110101",
38343 => "0000000001110101",38344 => "0000000001110101",
38345 => "0000000001110101",38346 => "0000000001110101",
38347 => "0000000001110101",38348 => "0000000001110101",
38349 => "0000000001110101",38350 => "0000000001110101",
38351 => "0000000001110101",38352 => "0000000001110101",
38353 => "0000000001110101",38354 => "0000000001110101",
38355 => "0000000001110101",38356 => "0000000001110101",
38357 => "0000000001110101",38358 => "0000000001110101",
38359 => "0000000001110101",38360 => "0000000001110101",
38361 => "0000000001110101",38362 => "0000000001110101",
38363 => "0000000001110100",38364 => "0000000001110100",
38365 => "0000000001110100",38366 => "0000000001110100",
38367 => "0000000001110100",38368 => "0000000001110100",
38369 => "0000000001110100",38370 => "0000000001110100",
38371 => "0000000001110100",38372 => "0000000001110100",
38373 => "0000000001110100",38374 => "0000000001110100",
38375 => "0000000001110100",38376 => "0000000001110100",
38377 => "0000000001110100",38378 => "0000000001110100",
38379 => "0000000001110100",38380 => "0000000001110100",
38381 => "0000000001110100",38382 => "0000000001110100",
38383 => "0000000001110100",38384 => "0000000001110100",
38385 => "0000000001110100",38386 => "0000000001110100",
38387 => "0000000001110100",38388 => "0000000001110100",
38389 => "0000000001110100",38390 => "0000000001110100",
38391 => "0000000001110100",38392 => "0000000001110100",
38393 => "0000000001110100",38394 => "0000000001110100",
38395 => "0000000001110100",38396 => "0000000001110100",
38397 => "0000000001110100",38398 => "0000000001110100",
38399 => "0000000001110100",38400 => "0000000001110100",
38401 => "0000000001110100",38402 => "0000000001110100",
38403 => "0000000001110100",38404 => "0000000001110100",
38405 => "0000000001110100",38406 => "0000000001110100",
38407 => "0000000001110100",38408 => "0000000001110100",
38409 => "0000000001110100",38410 => "0000000001110100",
38411 => "0000000001110100",38412 => "0000000001110100",
38413 => "0000000001110100",38414 => "0000000001110100",
38415 => "0000000001110100",38416 => "0000000001110100",
38417 => "0000000001110100",38418 => "0000000001110100",
38419 => "0000000001110100",38420 => "0000000001110100",
38421 => "0000000001110100",38422 => "0000000001110100",
38423 => "0000000001110100",38424 => "0000000001110100",
38425 => "0000000001110100",38426 => "0000000001110100",
38427 => "0000000001110100",38428 => "0000000001110100",
38429 => "0000000001110100",38430 => "0000000001110100",
38431 => "0000000001110100",38432 => "0000000001110100",
38433 => "0000000001110100",38434 => "0000000001110100",
38435 => "0000000001110100",38436 => "0000000001110100",
38437 => "0000000001110100",38438 => "0000000001110100",
38439 => "0000000001110100",38440 => "0000000001110100",
38441 => "0000000001110100",38442 => "0000000001110100",
38443 => "0000000001110100",38444 => "0000000001110100",
38445 => "0000000001110100",38446 => "0000000001110100",
38447 => "0000000001110100",38448 => "0000000001110100",
38449 => "0000000001110011",38450 => "0000000001110011",
38451 => "0000000001110011",38452 => "0000000001110011",
38453 => "0000000001110011",38454 => "0000000001110011",
38455 => "0000000001110011",38456 => "0000000001110011",
38457 => "0000000001110011",38458 => "0000000001110011",
38459 => "0000000001110011",38460 => "0000000001110011",
38461 => "0000000001110011",38462 => "0000000001110011",
38463 => "0000000001110011",38464 => "0000000001110011",
38465 => "0000000001110011",38466 => "0000000001110011",
38467 => "0000000001110011",38468 => "0000000001110011",
38469 => "0000000001110011",38470 => "0000000001110011",
38471 => "0000000001110011",38472 => "0000000001110011",
38473 => "0000000001110011",38474 => "0000000001110011",
38475 => "0000000001110011",38476 => "0000000001110011",
38477 => "0000000001110011",38478 => "0000000001110011",
38479 => "0000000001110011",38480 => "0000000001110011",
38481 => "0000000001110011",38482 => "0000000001110011",
38483 => "0000000001110011",38484 => "0000000001110011",
38485 => "0000000001110011",38486 => "0000000001110011",
38487 => "0000000001110011",38488 => "0000000001110011",
38489 => "0000000001110011",38490 => "0000000001110011",
38491 => "0000000001110011",38492 => "0000000001110011",
38493 => "0000000001110011",38494 => "0000000001110011",
38495 => "0000000001110011",38496 => "0000000001110011",
38497 => "0000000001110011",38498 => "0000000001110011",
38499 => "0000000001110011",38500 => "0000000001110011",
38501 => "0000000001110011",38502 => "0000000001110011",
38503 => "0000000001110011",38504 => "0000000001110011",
38505 => "0000000001110011",38506 => "0000000001110011",
38507 => "0000000001110011",38508 => "0000000001110011",
38509 => "0000000001110011",38510 => "0000000001110011",
38511 => "0000000001110011",38512 => "0000000001110011",
38513 => "0000000001110011",38514 => "0000000001110011",
38515 => "0000000001110011",38516 => "0000000001110011",
38517 => "0000000001110011",38518 => "0000000001110011",
38519 => "0000000001110011",38520 => "0000000001110011",
38521 => "0000000001110011",38522 => "0000000001110011",
38523 => "0000000001110011",38524 => "0000000001110011",
38525 => "0000000001110011",38526 => "0000000001110011",
38527 => "0000000001110011",38528 => "0000000001110011",
38529 => "0000000001110011",38530 => "0000000001110011",
38531 => "0000000001110011",38532 => "0000000001110011",
38533 => "0000000001110011",38534 => "0000000001110011",
38535 => "0000000001110011",38536 => "0000000001110010",
38537 => "0000000001110010",38538 => "0000000001110010",
38539 => "0000000001110010",38540 => "0000000001110010",
38541 => "0000000001110010",38542 => "0000000001110010",
38543 => "0000000001110010",38544 => "0000000001110010",
38545 => "0000000001110010",38546 => "0000000001110010",
38547 => "0000000001110010",38548 => "0000000001110010",
38549 => "0000000001110010",38550 => "0000000001110010",
38551 => "0000000001110010",38552 => "0000000001110010",
38553 => "0000000001110010",38554 => "0000000001110010",
38555 => "0000000001110010",38556 => "0000000001110010",
38557 => "0000000001110010",38558 => "0000000001110010",
38559 => "0000000001110010",38560 => "0000000001110010",
38561 => "0000000001110010",38562 => "0000000001110010",
38563 => "0000000001110010",38564 => "0000000001110010",
38565 => "0000000001110010",38566 => "0000000001110010",
38567 => "0000000001110010",38568 => "0000000001110010",
38569 => "0000000001110010",38570 => "0000000001110010",
38571 => "0000000001110010",38572 => "0000000001110010",
38573 => "0000000001110010",38574 => "0000000001110010",
38575 => "0000000001110010",38576 => "0000000001110010",
38577 => "0000000001110010",38578 => "0000000001110010",
38579 => "0000000001110010",38580 => "0000000001110010",
38581 => "0000000001110010",38582 => "0000000001110010",
38583 => "0000000001110010",38584 => "0000000001110010",
38585 => "0000000001110010",38586 => "0000000001110010",
38587 => "0000000001110010",38588 => "0000000001110010",
38589 => "0000000001110010",38590 => "0000000001110010",
38591 => "0000000001110010",38592 => "0000000001110010",
38593 => "0000000001110010",38594 => "0000000001110010",
38595 => "0000000001110010",38596 => "0000000001110010",
38597 => "0000000001110010",38598 => "0000000001110010",
38599 => "0000000001110010",38600 => "0000000001110010",
38601 => "0000000001110010",38602 => "0000000001110010",
38603 => "0000000001110010",38604 => "0000000001110010",
38605 => "0000000001110010",38606 => "0000000001110010",
38607 => "0000000001110010",38608 => "0000000001110010",
38609 => "0000000001110010",38610 => "0000000001110010",
38611 => "0000000001110010",38612 => "0000000001110010",
38613 => "0000000001110010",38614 => "0000000001110010",
38615 => "0000000001110010",38616 => "0000000001110010",
38617 => "0000000001110010",38618 => "0000000001110010",
38619 => "0000000001110010",38620 => "0000000001110010",
38621 => "0000000001110010",38622 => "0000000001110010",
38623 => "0000000001110010",38624 => "0000000001110001",
38625 => "0000000001110001",38626 => "0000000001110001",
38627 => "0000000001110001",38628 => "0000000001110001",
38629 => "0000000001110001",38630 => "0000000001110001",
38631 => "0000000001110001",38632 => "0000000001110001",
38633 => "0000000001110001",38634 => "0000000001110001",
38635 => "0000000001110001",38636 => "0000000001110001",
38637 => "0000000001110001",38638 => "0000000001110001",
38639 => "0000000001110001",38640 => "0000000001110001",
38641 => "0000000001110001",38642 => "0000000001110001",
38643 => "0000000001110001",38644 => "0000000001110001",
38645 => "0000000001110001",38646 => "0000000001110001",
38647 => "0000000001110001",38648 => "0000000001110001",
38649 => "0000000001110001",38650 => "0000000001110001",
38651 => "0000000001110001",38652 => "0000000001110001",
38653 => "0000000001110001",38654 => "0000000001110001",
38655 => "0000000001110001",38656 => "0000000001110001",
38657 => "0000000001110001",38658 => "0000000001110001",
38659 => "0000000001110001",38660 => "0000000001110001",
38661 => "0000000001110001",38662 => "0000000001110001",
38663 => "0000000001110001",38664 => "0000000001110001",
38665 => "0000000001110001",38666 => "0000000001110001",
38667 => "0000000001110001",38668 => "0000000001110001",
38669 => "0000000001110001",38670 => "0000000001110001",
38671 => "0000000001110001",38672 => "0000000001110001",
38673 => "0000000001110001",38674 => "0000000001110001",
38675 => "0000000001110001",38676 => "0000000001110001",
38677 => "0000000001110001",38678 => "0000000001110001",
38679 => "0000000001110001",38680 => "0000000001110001",
38681 => "0000000001110001",38682 => "0000000001110001",
38683 => "0000000001110001",38684 => "0000000001110001",
38685 => "0000000001110001",38686 => "0000000001110001",
38687 => "0000000001110001",38688 => "0000000001110001",
38689 => "0000000001110001",38690 => "0000000001110001",
38691 => "0000000001110001",38692 => "0000000001110001",
38693 => "0000000001110001",38694 => "0000000001110001",
38695 => "0000000001110001",38696 => "0000000001110001",
38697 => "0000000001110001",38698 => "0000000001110001",
38699 => "0000000001110001",38700 => "0000000001110001",
38701 => "0000000001110001",38702 => "0000000001110001",
38703 => "0000000001110001",38704 => "0000000001110001",
38705 => "0000000001110001",38706 => "0000000001110001",
38707 => "0000000001110001",38708 => "0000000001110001",
38709 => "0000000001110001",38710 => "0000000001110001",
38711 => "0000000001110001",38712 => "0000000001110001",
38713 => "0000000001110000",38714 => "0000000001110000",
38715 => "0000000001110000",38716 => "0000000001110000",
38717 => "0000000001110000",38718 => "0000000001110000",
38719 => "0000000001110000",38720 => "0000000001110000",
38721 => "0000000001110000",38722 => "0000000001110000",
38723 => "0000000001110000",38724 => "0000000001110000",
38725 => "0000000001110000",38726 => "0000000001110000",
38727 => "0000000001110000",38728 => "0000000001110000",
38729 => "0000000001110000",38730 => "0000000001110000",
38731 => "0000000001110000",38732 => "0000000001110000",
38733 => "0000000001110000",38734 => "0000000001110000",
38735 => "0000000001110000",38736 => "0000000001110000",
38737 => "0000000001110000",38738 => "0000000001110000",
38739 => "0000000001110000",38740 => "0000000001110000",
38741 => "0000000001110000",38742 => "0000000001110000",
38743 => "0000000001110000",38744 => "0000000001110000",
38745 => "0000000001110000",38746 => "0000000001110000",
38747 => "0000000001110000",38748 => "0000000001110000",
38749 => "0000000001110000",38750 => "0000000001110000",
38751 => "0000000001110000",38752 => "0000000001110000",
38753 => "0000000001110000",38754 => "0000000001110000",
38755 => "0000000001110000",38756 => "0000000001110000",
38757 => "0000000001110000",38758 => "0000000001110000",
38759 => "0000000001110000",38760 => "0000000001110000",
38761 => "0000000001110000",38762 => "0000000001110000",
38763 => "0000000001110000",38764 => "0000000001110000",
38765 => "0000000001110000",38766 => "0000000001110000",
38767 => "0000000001110000",38768 => "0000000001110000",
38769 => "0000000001110000",38770 => "0000000001110000",
38771 => "0000000001110000",38772 => "0000000001110000",
38773 => "0000000001110000",38774 => "0000000001110000",
38775 => "0000000001110000",38776 => "0000000001110000",
38777 => "0000000001110000",38778 => "0000000001110000",
38779 => "0000000001110000",38780 => "0000000001110000",
38781 => "0000000001110000",38782 => "0000000001110000",
38783 => "0000000001110000",38784 => "0000000001110000",
38785 => "0000000001110000",38786 => "0000000001110000",
38787 => "0000000001110000",38788 => "0000000001110000",
38789 => "0000000001110000",38790 => "0000000001110000",
38791 => "0000000001110000",38792 => "0000000001110000",
38793 => "0000000001110000",38794 => "0000000001110000",
38795 => "0000000001110000",38796 => "0000000001110000",
38797 => "0000000001110000",38798 => "0000000001110000",
38799 => "0000000001110000",38800 => "0000000001110000",
38801 => "0000000001110000",38802 => "0000000001101111",
38803 => "0000000001101111",38804 => "0000000001101111",
38805 => "0000000001101111",38806 => "0000000001101111",
38807 => "0000000001101111",38808 => "0000000001101111",
38809 => "0000000001101111",38810 => "0000000001101111",
38811 => "0000000001101111",38812 => "0000000001101111",
38813 => "0000000001101111",38814 => "0000000001101111",
38815 => "0000000001101111",38816 => "0000000001101111",
38817 => "0000000001101111",38818 => "0000000001101111",
38819 => "0000000001101111",38820 => "0000000001101111",
38821 => "0000000001101111",38822 => "0000000001101111",
38823 => "0000000001101111",38824 => "0000000001101111",
38825 => "0000000001101111",38826 => "0000000001101111",
38827 => "0000000001101111",38828 => "0000000001101111",
38829 => "0000000001101111",38830 => "0000000001101111",
38831 => "0000000001101111",38832 => "0000000001101111",
38833 => "0000000001101111",38834 => "0000000001101111",
38835 => "0000000001101111",38836 => "0000000001101111",
38837 => "0000000001101111",38838 => "0000000001101111",
38839 => "0000000001101111",38840 => "0000000001101111",
38841 => "0000000001101111",38842 => "0000000001101111",
38843 => "0000000001101111",38844 => "0000000001101111",
38845 => "0000000001101111",38846 => "0000000001101111",
38847 => "0000000001101111",38848 => "0000000001101111",
38849 => "0000000001101111",38850 => "0000000001101111",
38851 => "0000000001101111",38852 => "0000000001101111",
38853 => "0000000001101111",38854 => "0000000001101111",
38855 => "0000000001101111",38856 => "0000000001101111",
38857 => "0000000001101111",38858 => "0000000001101111",
38859 => "0000000001101111",38860 => "0000000001101111",
38861 => "0000000001101111",38862 => "0000000001101111",
38863 => "0000000001101111",38864 => "0000000001101111",
38865 => "0000000001101111",38866 => "0000000001101111",
38867 => "0000000001101111",38868 => "0000000001101111",
38869 => "0000000001101111",38870 => "0000000001101111",
38871 => "0000000001101111",38872 => "0000000001101111",
38873 => "0000000001101111",38874 => "0000000001101111",
38875 => "0000000001101111",38876 => "0000000001101111",
38877 => "0000000001101111",38878 => "0000000001101111",
38879 => "0000000001101111",38880 => "0000000001101111",
38881 => "0000000001101111",38882 => "0000000001101111",
38883 => "0000000001101111",38884 => "0000000001101111",
38885 => "0000000001101111",38886 => "0000000001101111",
38887 => "0000000001101111",38888 => "0000000001101111",
38889 => "0000000001101111",38890 => "0000000001101111",
38891 => "0000000001101111",38892 => "0000000000001011",
38893 => "0000000000001011",38894 => "0000000000001011",
38895 => "0000000000001011",38896 => "0000000000001011",
38897 => "0000000000001011",38898 => "0000000000001011",
38899 => "0000000000001011",38900 => "0000000000001011",
38901 => "0000000000001011",38902 => "0000000000001011",
38903 => "0000000000001011",38904 => "0000000000001011",
38905 => "0000000000001011",38906 => "0000000000001011",
38907 => "0000000000001011",38908 => "0000000000001011",
38909 => "0000000000001011",38910 => "0000000000001011",
38911 => "0000000000001011",38912 => "0000000000000101",
38913 => "0000000000101101",38914 => "0000000000101001",
38915 => "0000000000100101",38916 => "0000000000100001",
38917 => "0000000000000011",38918 => "0000000000011011",
38919 => "0000000000011001",38920 => "0000000000010110",
38921 => "0000000000000010",38922 => "0000000000101101",
38923 => "0000000000101101",38924 => "0000000000101100",
38925 => "0000000000101100",38926 => "0000000000101011",
38927 => "0000000000101011",38928 => "0000000000101010",
38929 => "0000000000101010",38930 => "0000000000101010",
38931 => "0000000000101001",38932 => "0000000000101001",
38933 => "0000000000000100",38934 => "0000000000000100",
38935 => "0000000000000100",38936 => "0000000000100111",
38937 => "0000000000100111",38938 => "0000000000100110",
38939 => "0000000000100110",38940 => "0000000000100110",
38941 => "0000000000100101",38942 => "0000000000100101",
38943 => "0000000000100101",38944 => "0000000000100100",
38945 => "0000000000100100",38946 => "0000000000100011",
38947 => "0000000000100011",38948 => "0000000000100011",
38949 => "0000000000100010",38950 => "0000000000100010",
38951 => "0000000000100010",38952 => "0000000000100001",
38953 => "0000000000100001",38954 => "0000000000100001",
38955 => "0000000000100000",38956 => "0000000000100000",
38957 => "0000000000100000",38958 => "0000000000011111",
38959 => "0000000000011111",38960 => "0000000000011111",
38961 => "0000000000011111",38962 => "0000000000000011",
38963 => "0000000000000011",38964 => "0000000000000011",
38965 => "0000000000011101",38966 => "0000000000011101",
38967 => "0000000000011101",38968 => "0000000000011100",
38969 => "0000000000011100",38970 => "0000000000011100",
38971 => "0000000000011100",38972 => "0000000000011011",
38973 => "0000000000011011",38974 => "0000000000011011",
38975 => "0000000000011011",38976 => "0000000000011010",
38977 => "0000000000011010",38978 => "0000000000011010",
38979 => "0000000000011001",38980 => "0000000000011001",
38981 => "0000000000011001",38982 => "0000000000011001",
38983 => "0000000000011000",38984 => "0000000000011000",
38985 => "0000000000011000",38986 => "0000000000011000",
38987 => "0000000000011000",38988 => "0000000000010111",
38989 => "0000000000010111",38990 => "0000000000010111",
38991 => "0000000000010111",38992 => "0000000000010110",
38993 => "0000000000010110",38994 => "0000000000010110",
38995 => "0000000000010110",38996 => "0000000000010101",
38997 => "0000000000010101",38998 => "0000000000010101",
38999 => "0000000000010101",39000 => "0000000000010101",
39001 => "0000000000000010",39002 => "0000000000000010",
39003 => "0000000000000010",39004 => "0000000000000010",
39005 => "0000000000000010",39006 => "0000000000010011",
39007 => "0000000000010011",39008 => "0000000000010011",
39009 => "0000000000010011",39010 => "0000000000010011",
39011 => "0000000000010010",39012 => "0000000000101101",
39013 => "0000000000101101",39014 => "0000000000101101",
39015 => "0000000000101101",39016 => "0000000000101101",
39017 => "0000000000101101",39018 => "0000000000101101",
39019 => "0000000000101101",39020 => "0000000000101101",
39021 => "0000000000101101",39022 => "0000000000101101",
39023 => "0000000000101101",39024 => "0000000000101101",
39025 => "0000000000101100",39026 => "0000000000101100",
39027 => "0000000000101100",39028 => "0000000000101100",
39029 => "0000000000101100",39030 => "0000000000101100",
39031 => "0000000000101100",39032 => "0000000000101100",
39033 => "0000000000101100",39034 => "0000000000101100",
39035 => "0000000000101100",39036 => "0000000000101100",
39037 => "0000000000101100",39038 => "0000000000101100",
39039 => "0000000000101100",39040 => "0000000000101100",
39041 => "0000000000101100",39042 => "0000000000101100",
39043 => "0000000000101100",39044 => "0000000000101100",
39045 => "0000000000101100",39046 => "0000000000101100",
39047 => "0000000000101011",39048 => "0000000000101011",
39049 => "0000000000101011",39050 => "0000000000101011",
39051 => "0000000000101011",39052 => "0000000000101011",
39053 => "0000000000101011",39054 => "0000000000101011",
39055 => "0000000000101011",39056 => "0000000000101011",
39057 => "0000000000101011",39058 => "0000000000101011",
39059 => "0000000000101011",39060 => "0000000000101011",
39061 => "0000000000101011",39062 => "0000000000101011",
39063 => "0000000000101011",39064 => "0000000000101011",
39065 => "0000000000101011",39066 => "0000000000101011",
39067 => "0000000000101011",39068 => "0000000000101011",
39069 => "0000000000101011",39070 => "0000000000101011",
39071 => "0000000000101010",39072 => "0000000000101010",
39073 => "0000000000101010",39074 => "0000000000101010",
39075 => "0000000000101010",39076 => "0000000000101010",
39077 => "0000000000101010",39078 => "0000000000101010",
39079 => "0000000000101010",39080 => "0000000000101010",
39081 => "0000000000101010",39082 => "0000000000101010",
39083 => "0000000000101010",39084 => "0000000000101010",
39085 => "0000000000101010",39086 => "0000000000101010",
39087 => "0000000000101010",39088 => "0000000000101010",
39089 => "0000000000101010",39090 => "0000000000101010",
39091 => "0000000000101010",39092 => "0000000000101010",
39093 => "0000000000101010",39094 => "0000000000101010",
39095 => "0000000000101001",39096 => "0000000000101001",
39097 => "0000000000101001",39098 => "0000000000101001",
39099 => "0000000000101001",39100 => "0000000000101001",
39101 => "0000000000101001",39102 => "0000000000101001",
39103 => "0000000000101001",39104 => "0000000000101001",
39105 => "0000000000101001",39106 => "0000000000101001",
39107 => "0000000000101001",39108 => "0000000000101001",
39109 => "0000000000101001",39110 => "0000000000101001",
39111 => "0000000000101001",39112 => "0000000000101001",
39113 => "0000000000101001",39114 => "0000000000101001",
39115 => "0000000000101001",39116 => "0000000000101001",
39117 => "0000000000101001",39118 => "0000000000101001",
39119 => "0000000000000100",39120 => "0000000000000100",
39121 => "0000000000000100",39122 => "0000000000000100",
39123 => "0000000000000100",39124 => "0000000000000100",
39125 => "0000000000000100",39126 => "0000000000000100",
39127 => "0000000000000100",39128 => "0000000000000100",
39129 => "0000000000000100",39130 => "0000000000000100",
39131 => "0000000000000100",39132 => "0000000000000100",
39133 => "0000000000000100",39134 => "0000000000000100",
39135 => "0000000000000100",39136 => "0000000000000100",
39137 => "0000000000000100",39138 => "0000000000000100",
39139 => "0000000000000100",39140 => "0000000000000100",
39141 => "0000000000000100",39142 => "0000000000000100",
39143 => "0000000000000100",39144 => "0000000000100111",
39145 => "0000000000100111",39146 => "0000000000100111",
39147 => "0000000000100111",39148 => "0000000000100111",
39149 => "0000000000100111",39150 => "0000000000100111",
39151 => "0000000000100111",39152 => "0000000000100111",
39153 => "0000000000100111",39154 => "0000000000100111",
39155 => "0000000000100111",39156 => "0000000000100111",
39157 => "0000000000100111",39158 => "0000000000100111",
39159 => "0000000000100111",39160 => "0000000000100111",
39161 => "0000000000100111",39162 => "0000000000100111",
39163 => "0000000000100111",39164 => "0000000000100111",
39165 => "0000000000100111",39166 => "0000000000100111",
39167 => "0000000000100111",39168 => "0000000000100111",
39169 => "0000000000100111",39170 => "0000000000100110",
39171 => "0000000000100110",39172 => "0000000000100110",
39173 => "0000000000100110",39174 => "0000000000100110",
39175 => "0000000000100110",39176 => "0000000000100110",
39177 => "0000000000100110",39178 => "0000000000100110",
39179 => "0000000000100110",39180 => "0000000000100110",
39181 => "0000000000100110",39182 => "0000000000100110",
39183 => "0000000000100110",39184 => "0000000000100110",
39185 => "0000000000100110",39186 => "0000000000100110",
39187 => "0000000000100110",39188 => "0000000000100110",
39189 => "0000000000100110",39190 => "0000000000100110",
39191 => "0000000000100110",39192 => "0000000000100110",
39193 => "0000000000100110",39194 => "0000000000100110",
39195 => "0000000000100110",39196 => "0000000000100101",
39197 => "0000000000100101",39198 => "0000000000100101",
39199 => "0000000000100101",39200 => "0000000000100101",
39201 => "0000000000100101",39202 => "0000000000100101",
39203 => "0000000000100101",39204 => "0000000000100101",
39205 => "0000000000100101",39206 => "0000000000100101",
39207 => "0000000000100101",39208 => "0000000000100101",
39209 => "0000000000100101",39210 => "0000000000100101",
39211 => "0000000000100101",39212 => "0000000000100101",
39213 => "0000000000100101",39214 => "0000000000100101",
39215 => "0000000000100101",39216 => "0000000000100101",
39217 => "0000000000100101",39218 => "0000000000100101",
39219 => "0000000000100101",39220 => "0000000000100101",
39221 => "0000000000100101",39222 => "0000000000100101",
39223 => "0000000000100100",39224 => "0000000000100100",
39225 => "0000000000100100",39226 => "0000000000100100",
39227 => "0000000000100100",39228 => "0000000000100100",
39229 => "0000000000100100",39230 => "0000000000100100",
39231 => "0000000000100100",39232 => "0000000000100100",
39233 => "0000000000100100",39234 => "0000000000100100",
39235 => "0000000000100100",39236 => "0000000000100100",
39237 => "0000000000100100",39238 => "0000000000100100",
39239 => "0000000000100100",39240 => "0000000000100100",
39241 => "0000000000100100",39242 => "0000000000100100",
39243 => "0000000000100100",39244 => "0000000000100100",
39245 => "0000000000100100",39246 => "0000000000100100",
39247 => "0000000000100100",39248 => "0000000000100100",
39249 => "0000000000100100",39250 => "0000000000100100",
39251 => "0000000000100011",39252 => "0000000000100011",
39253 => "0000000000100011",39254 => "0000000000100011",
39255 => "0000000000100011",39256 => "0000000000100011",
39257 => "0000000000100011",39258 => "0000000000100011",
39259 => "0000000000100011",39260 => "0000000000100011",
39261 => "0000000000100011",39262 => "0000000000100011",
39263 => "0000000000100011",39264 => "0000000000100011",
39265 => "0000000000100011",39266 => "0000000000100011",
39267 => "0000000000100011",39268 => "0000000000100011",
39269 => "0000000000100011",39270 => "0000000000100011",
39271 => "0000000000100011",39272 => "0000000000100011",
39273 => "0000000000100011",39274 => "0000000000100011",
39275 => "0000000000100011",39276 => "0000000000100011",
39277 => "0000000000100011",39278 => "0000000000100011",
39279 => "0000000000100010",39280 => "0000000000100010",
39281 => "0000000000100010",39282 => "0000000000100010",
39283 => "0000000000100010",39284 => "0000000000100010",
39285 => "0000000000100010",39286 => "0000000000100010",
39287 => "0000000000100010",39288 => "0000000000100010",
39289 => "0000000000100010",39290 => "0000000000100010",
39291 => "0000000000100010",39292 => "0000000000100010",
39293 => "0000000000100010",39294 => "0000000000100010",
39295 => "0000000000100010",39296 => "0000000000100010",
39297 => "0000000000100010",39298 => "0000000000100010",
39299 => "0000000000100010",39300 => "0000000000100010",
39301 => "0000000000100010",39302 => "0000000000100010",
39303 => "0000000000100010",39304 => "0000000000100010",
39305 => "0000000000100010",39306 => "0000000000100010",
39307 => "0000000000100010",39308 => "0000000000100010",
39309 => "0000000000100001",39310 => "0000000000100001",
39311 => "0000000000100001",39312 => "0000000000100001",
39313 => "0000000000100001",39314 => "0000000000100001",
39315 => "0000000000100001",39316 => "0000000000100001",
39317 => "0000000000100001",39318 => "0000000000100001",
39319 => "0000000000100001",39320 => "0000000000100001",
39321 => "0000000000100001",39322 => "0000000000100001",
39323 => "0000000000100001",39324 => "0000000000100001",
39325 => "0000000000100001",39326 => "0000000000100001",
39327 => "0000000000100001",39328 => "0000000000100001",
39329 => "0000000000100001",39330 => "0000000000100001",
39331 => "0000000000100001",39332 => "0000000000100001",
39333 => "0000000000100001",39334 => "0000000000100001",
39335 => "0000000000100001",39336 => "0000000000100001",
39337 => "0000000000100001",39338 => "0000000000100001",
39339 => "0000000000100000",39340 => "0000000000100000",
39341 => "0000000000100000",39342 => "0000000000100000",
39343 => "0000000000100000",39344 => "0000000000100000",
39345 => "0000000000100000",39346 => "0000000000100000",
39347 => "0000000000100000",39348 => "0000000000100000",
39349 => "0000000000100000",39350 => "0000000000100000",
39351 => "0000000000100000",39352 => "0000000000100000",
39353 => "0000000000100000",39354 => "0000000000100000",
39355 => "0000000000100000",39356 => "0000000000100000",
39357 => "0000000000100000",39358 => "0000000000100000",
39359 => "0000000000100000",39360 => "0000000000100000",
39361 => "0000000000100000",39362 => "0000000000100000",
39363 => "0000000000100000",39364 => "0000000000100000",
39365 => "0000000000100000",39366 => "0000000000100000",
39367 => "0000000000100000",39368 => "0000000000100000",
39369 => "0000000000100000",39370 => "0000000000011111",
39371 => "0000000000011111",39372 => "0000000000011111",
39373 => "0000000000011111",39374 => "0000000000011111",
39375 => "0000000000011111",39376 => "0000000000011111",
39377 => "0000000000011111",39378 => "0000000000011111",
39379 => "0000000000011111",39380 => "0000000000011111",
39381 => "0000000000011111",39382 => "0000000000011111",
39383 => "0000000000011111",39384 => "0000000000011111",
39385 => "0000000000011111",39386 => "0000000000011111",
39387 => "0000000000011111",39388 => "0000000000011111",
39389 => "0000000000011111",39390 => "0000000000011111",
39391 => "0000000000011111",39392 => "0000000000011111",
39393 => "0000000000011111",39394 => "0000000000011111",
39395 => "0000000000011111",39396 => "0000000000011111",
39397 => "0000000000011111",39398 => "0000000000011111",
39399 => "0000000000011111",39400 => "0000000000011111",
39401 => "0000000000011111",39402 => "0000000000011111",
39403 => "0000000000000011",39404 => "0000000000000011",
39405 => "0000000000000011",39406 => "0000000000000011",
39407 => "0000000000000011",39408 => "0000000000000011",
39409 => "0000000000000011",39410 => "0000000000000011",
39411 => "0000000000000011",39412 => "0000000000000011",
39413 => "0000000000000011",39414 => "0000000000000011",
39415 => "0000000000000011",39416 => "0000000000000011",
39417 => "0000000000000011",39418 => "0000000000000011",
39419 => "0000000000000011",39420 => "0000000000000011",
39421 => "0000000000000011",39422 => "0000000000000011",
39423 => "0000000000000011",39424 => "0000000000000011",
39425 => "0000000000000011",39426 => "0000000000000011",
39427 => "0000000000000011",39428 => "0000000000000011",
39429 => "0000000000000011",39430 => "0000000000000011",
39431 => "0000000000000011",39432 => "0000000000000011",
39433 => "0000000000000011",39434 => "0000000000000011",
39435 => "0000000000000011",39436 => "0000000000011101",
39437 => "0000000000011101",39438 => "0000000000011101",
39439 => "0000000000011101",39440 => "0000000000011101",
39441 => "0000000000011101",39442 => "0000000000011101",
39443 => "0000000000011101",39444 => "0000000000011101",
39445 => "0000000000011101",39446 => "0000000000011101",
39447 => "0000000000011101",39448 => "0000000000011101",
39449 => "0000000000011101",39450 => "0000000000011101",
39451 => "0000000000011101",39452 => "0000000000011101",
39453 => "0000000000011101",39454 => "0000000000011101",
39455 => "0000000000011101",39456 => "0000000000011101",
39457 => "0000000000011101",39458 => "0000000000011101",
39459 => "0000000000011101",39460 => "0000000000011101",
39461 => "0000000000011101",39462 => "0000000000011101",
39463 => "0000000000011101",39464 => "0000000000011101",
39465 => "0000000000011101",39466 => "0000000000011101",
39467 => "0000000000011101",39468 => "0000000000011101",
39469 => "0000000000011101",39470 => "0000000000011100",
39471 => "0000000000011100",39472 => "0000000000011100",
39473 => "0000000000011100",39474 => "0000000000011100",
39475 => "0000000000011100",39476 => "0000000000011100",
39477 => "0000000000011100",39478 => "0000000000011100",
39479 => "0000000000011100",39480 => "0000000000011100",
39481 => "0000000000011100",39482 => "0000000000011100",
39483 => "0000000000011100",39484 => "0000000000011100",
39485 => "0000000000011100",39486 => "0000000000011100",
39487 => "0000000000011100",39488 => "0000000000011100",
39489 => "0000000000011100",39490 => "0000000000011100",
39491 => "0000000000011100",39492 => "0000000000011100",
39493 => "0000000000011100",39494 => "0000000000011100",
39495 => "0000000000011100",39496 => "0000000000011100",
39497 => "0000000000011100",39498 => "0000000000011100",
39499 => "0000000000011100",39500 => "0000000000011100",
39501 => "0000000000011100",39502 => "0000000000011100",
39503 => "0000000000011100",39504 => "0000000000011100",
39505 => "0000000000011100",39506 => "0000000000011011",
39507 => "0000000000011011",39508 => "0000000000011011",
39509 => "0000000000011011",39510 => "0000000000011011",
39511 => "0000000000011011",39512 => "0000000000011011",
39513 => "0000000000011011",39514 => "0000000000011011",
39515 => "0000000000011011",39516 => "0000000000011011",
39517 => "0000000000011011",39518 => "0000000000011011",
39519 => "0000000000011011",39520 => "0000000000011011",
39521 => "0000000000011011",39522 => "0000000000011011",
39523 => "0000000000011011",39524 => "0000000000011011",
39525 => "0000000000011011",39526 => "0000000000011011",
39527 => "0000000000011011",39528 => "0000000000011011",
39529 => "0000000000011011",39530 => "0000000000011011",
39531 => "0000000000011011",39532 => "0000000000011011",
39533 => "0000000000011011",39534 => "0000000000011011",
39535 => "0000000000011011",39536 => "0000000000011011",
39537 => "0000000000011011",39538 => "0000000000011011",
39539 => "0000000000011011",39540 => "0000000000011011",
39541 => "0000000000011011",39542 => "0000000000011011",
39543 => "0000000000011010",39544 => "0000000000011010",
39545 => "0000000000011010",39546 => "0000000000011010",
39547 => "0000000000011010",39548 => "0000000000011010",
39549 => "0000000000011010",39550 => "0000000000011010",
39551 => "0000000000011010",39552 => "0000000000011010",
39553 => "0000000000011010",39554 => "0000000000011010",
39555 => "0000000000011010",39556 => "0000000000011010",
39557 => "0000000000011010",39558 => "0000000000011010",
39559 => "0000000000011010",39560 => "0000000000011010",
39561 => "0000000000011010",39562 => "0000000000011010",
39563 => "0000000000011010",39564 => "0000000000011010",
39565 => "0000000000011010",39566 => "0000000000011010",
39567 => "0000000000011010",39568 => "0000000000011010",
39569 => "0000000000011010",39570 => "0000000000011010",
39571 => "0000000000011010",39572 => "0000000000011010",
39573 => "0000000000011010",39574 => "0000000000011010",
39575 => "0000000000011010",39576 => "0000000000011010",
39577 => "0000000000011010",39578 => "0000000000011010",
39579 => "0000000000011010",39580 => "0000000000011010",
39581 => "0000000000011010",39582 => "0000000000011001",
39583 => "0000000000011001",39584 => "0000000000011001",
39585 => "0000000000011001",39586 => "0000000000011001",
39587 => "0000000000011001",39588 => "0000000000011001",
39589 => "0000000000011001",39590 => "0000000000011001",
39591 => "0000000000011001",39592 => "0000000000011001",
39593 => "0000000000011001",39594 => "0000000000011001",
39595 => "0000000000011001",39596 => "0000000000011001",
39597 => "0000000000011001",39598 => "0000000000011001",
39599 => "0000000000011001",39600 => "0000000000011001",
39601 => "0000000000011001",39602 => "0000000000011001",
39603 => "0000000000011001",39604 => "0000000000011001",
39605 => "0000000000011001",39606 => "0000000000011001",
39607 => "0000000000011001",39608 => "0000000000011001",
39609 => "0000000000011001",39610 => "0000000000011001",
39611 => "0000000000011001",39612 => "0000000000011001",
39613 => "0000000000011001",39614 => "0000000000011001",
39615 => "0000000000011001",39616 => "0000000000011001",
39617 => "0000000000011001",39618 => "0000000000011001",
39619 => "0000000000011001",39620 => "0000000000011001",
39621 => "0000000000011001",39622 => "0000000000011000",
39623 => "0000000000011000",39624 => "0000000000011000",
39625 => "0000000000011000",39626 => "0000000000011000",
39627 => "0000000000011000",39628 => "0000000000011000",
39629 => "0000000000011000",39630 => "0000000000011000",
39631 => "0000000000011000",39632 => "0000000000011000",
39633 => "0000000000011000",39634 => "0000000000011000",
39635 => "0000000000011000",39636 => "0000000000011000",
39637 => "0000000000011000",39638 => "0000000000011000",
39639 => "0000000000011000",39640 => "0000000000011000",
39641 => "0000000000011000",39642 => "0000000000011000",
39643 => "0000000000011000",39644 => "0000000000011000",
39645 => "0000000000011000",39646 => "0000000000011000",
39647 => "0000000000011000",39648 => "0000000000011000",
39649 => "0000000000011000",39650 => "0000000000011000",
39651 => "0000000000011000",39652 => "0000000000011000",
39653 => "0000000000011000",39654 => "0000000000011000",
39655 => "0000000000011000",39656 => "0000000000011000",
39657 => "0000000000011000",39658 => "0000000000011000",
39659 => "0000000000011000",39660 => "0000000000011000",
39661 => "0000000000011000",39662 => "0000000000011000",
39663 => "0000000000010111",39664 => "0000000000010111",
39665 => "0000000000010111",39666 => "0000000000010111",
39667 => "0000000000010111",39668 => "0000000000010111",
39669 => "0000000000010111",39670 => "0000000000010111",
39671 => "0000000000010111",39672 => "0000000000010111",
39673 => "0000000000010111",39674 => "0000000000010111",
39675 => "0000000000010111",39676 => "0000000000010111",
39677 => "0000000000010111",39678 => "0000000000010111",
39679 => "0000000000010111",39680 => "0000000000010111",
39681 => "0000000000010111",39682 => "0000000000010111",
39683 => "0000000000010111",39684 => "0000000000010111",
39685 => "0000000000010111",39686 => "0000000000010111",
39687 => "0000000000010111",39688 => "0000000000010111",
39689 => "0000000000010111",39690 => "0000000000010111",
39691 => "0000000000010111",39692 => "0000000000010111",
39693 => "0000000000010111",39694 => "0000000000010111",
39695 => "0000000000010111",39696 => "0000000000010111",
39697 => "0000000000010111",39698 => "0000000000010111",
39699 => "0000000000010111",39700 => "0000000000010111",
39701 => "0000000000010111",39702 => "0000000000010111",
39703 => "0000000000010111",39704 => "0000000000010111",
39705 => "0000000000010111",39706 => "0000000000010111",
39707 => "0000000000010110",39708 => "0000000000010110",
39709 => "0000000000010110",39710 => "0000000000010110",
39711 => "0000000000010110",39712 => "0000000000010110",
39713 => "0000000000010110",39714 => "0000000000010110",
39715 => "0000000000010110",39716 => "0000000000010110",
39717 => "0000000000010110",39718 => "0000000000010110",
39719 => "0000000000010110",39720 => "0000000000010110",
39721 => "0000000000010110",39722 => "0000000000010110",
39723 => "0000000000010110",39724 => "0000000000010110",
39725 => "0000000000010110",39726 => "0000000000010110",
39727 => "0000000000010110",39728 => "0000000000010110",
39729 => "0000000000010110",39730 => "0000000000010110",
39731 => "0000000000010110",39732 => "0000000000010110",
39733 => "0000000000010110",39734 => "0000000000010110",
39735 => "0000000000010110",39736 => "0000000000010110",
39737 => "0000000000010110",39738 => "0000000000010110",
39739 => "0000000000010110",39740 => "0000000000010110",
39741 => "0000000000010110",39742 => "0000000000010110",
39743 => "0000000000010110",39744 => "0000000000010110",
39745 => "0000000000010110",39746 => "0000000000010110",
39747 => "0000000000010110",39748 => "0000000000010110",
39749 => "0000000000010110",39750 => "0000000000010110",
39751 => "0000000000010110",39752 => "0000000000010101",
39753 => "0000000000010101",39754 => "0000000000010101",
39755 => "0000000000010101",39756 => "0000000000010101",
39757 => "0000000000010101",39758 => "0000000000010101",
39759 => "0000000000010101",39760 => "0000000000010101",
39761 => "0000000000010101",39762 => "0000000000010101",
39763 => "0000000000010101",39764 => "0000000000010101",
39765 => "0000000000010101",39766 => "0000000000010101",
39767 => "0000000000010101",39768 => "0000000000010101",
39769 => "0000000000010101",39770 => "0000000000010101",
39771 => "0000000000010101",39772 => "0000000000010101",
39773 => "0000000000010101",39774 => "0000000000010101",
39775 => "0000000000010101",39776 => "0000000000010101",
39777 => "0000000000010101",39778 => "0000000000010101",
39779 => "0000000000010101",39780 => "0000000000010101",
39781 => "0000000000010101",39782 => "0000000000010101",
39783 => "0000000000010101",39784 => "0000000000010101",
39785 => "0000000000010101",39786 => "0000000000010101",
39787 => "0000000000010101",39788 => "0000000000010101",
39789 => "0000000000010101",39790 => "0000000000010101",
39791 => "0000000000010101",39792 => "0000000000010101",
39793 => "0000000000010101",39794 => "0000000000010101",
39795 => "0000000000010101",39796 => "0000000000010101",
39797 => "0000000000010101",39798 => "0000000000010101",
39799 => "0000000000010101",39800 => "0000000000000010",
39801 => "0000000000000010",39802 => "0000000000000010",
39803 => "0000000000000010",39804 => "0000000000000010",
39805 => "0000000000000010",39806 => "0000000000000010",
39807 => "0000000000000010",39808 => "0000000000000010",
39809 => "0000000000000010",39810 => "0000000000000010",
39811 => "0000000000000010",39812 => "0000000000000010",
39813 => "0000000000000010",39814 => "0000000000000010",
39815 => "0000000000000010",39816 => "0000000000000010",
39817 => "0000000000000010",39818 => "0000000000000010",
39819 => "0000000000000010",39820 => "0000000000000010",
39821 => "0000000000000010",39822 => "0000000000000010",
39823 => "0000000000000010",39824 => "0000000000000010",
39825 => "0000000000000010",39826 => "0000000000000010",
39827 => "0000000000000010",39828 => "0000000000000010",
39829 => "0000000000000010",39830 => "0000000000000010",
39831 => "0000000000000010",39832 => "0000000000000010",
39833 => "0000000000000010",39834 => "0000000000000010",
39835 => "0000000000000010",39836 => "0000000000000010",
39837 => "0000000000000010",39838 => "0000000000000010",
39839 => "0000000000000010",39840 => "0000000000000010",
39841 => "0000000000000010",39842 => "0000000000000010",
39843 => "0000000000000010",39844 => "0000000000000010",
39845 => "0000000000000010",39846 => "0000000000000010",
39847 => "0000000000000010",39848 => "0000000000000010",
39849 => "0000000000000010",39850 => "0000000000010011",
39851 => "0000000000010011",39852 => "0000000000010011",
39853 => "0000000000010011",39854 => "0000000000010011",
39855 => "0000000000010011",39856 => "0000000000010011",
39857 => "0000000000010011",39858 => "0000000000010011",
39859 => "0000000000010011",39860 => "0000000000010011",
39861 => "0000000000010011",39862 => "0000000000010011",
39863 => "0000000000010011",39864 => "0000000000010011",
39865 => "0000000000010011",39866 => "0000000000010011",
39867 => "0000000000010011",39868 => "0000000000010011",
39869 => "0000000000010011",39870 => "0000000000010011",
39871 => "0000000000010011",39872 => "0000000000010011",
39873 => "0000000000010011",39874 => "0000000000010011",
39875 => "0000000000010011",39876 => "0000000000010011",
39877 => "0000000000010011",39878 => "0000000000010011",
39879 => "0000000000010011",39880 => "0000000000010011",
39881 => "0000000000010011",39882 => "0000000000010011",
39883 => "0000000000010011",39884 => "0000000000010011",
39885 => "0000000000010011",39886 => "0000000000010011",
39887 => "0000000000010011",39888 => "0000000000010011",
39889 => "0000000000010011",39890 => "0000000000010011",
39891 => "0000000000010011",39892 => "0000000000010011",
39893 => "0000000000010011",39894 => "0000000000010011",
39895 => "0000000000010011",39896 => "0000000000010011",
39897 => "0000000000010011",39898 => "0000000000010011",
39899 => "0000000000010011",39900 => "0000000000010011",
39901 => "0000000000010011",39902 => "0000000000010010",
39903 => "0000000000010010",39904 => "0000000000010010",
39905 => "0000000000010010",39906 => "0000000000010010",
39907 => "0000000000010010",39908 => "0000000000010010",
39909 => "0000000000010010",39910 => "0000000000010010",
39911 => "0000000000010010",39912 => "0000000000101101",
39913 => "0000000000101101",39914 => "0000000000101101",
39915 => "0000000000101101",39916 => "0000000000101101",
39917 => "0000000000101101",39918 => "0000000000101101",
39919 => "0000000000101101",39920 => "0000000000101101",
39921 => "0000000000101101",39922 => "0000000000101101",
39923 => "0000000000101101",39924 => "0000000000101101",
39925 => "0000000000101101",39926 => "0000000000101101",
39927 => "0000000000101101",39928 => "0000000000101101",
39929 => "0000000000101101",39930 => "0000000000101101",
39931 => "0000000000101101",39932 => "0000000000101101",
39933 => "0000000000101101",39934 => "0000000000101101",
39935 => "0000000000101101",39936 => "0000000000101101",
39937 => "0000000000101101",39938 => "0000000000101101",
39939 => "0000000000101101",39940 => "0000000000101101",
39941 => "0000000000101101",39942 => "0000000000101101",
39943 => "0000000000101101",39944 => "0000000000101101",
39945 => "0000000000101101",39946 => "0000000000101101",
39947 => "0000000000101101",39948 => "0000000000101101",
39949 => "0000000000101101",39950 => "0000000000101101",
39951 => "0000000000101101",39952 => "0000000000101101",
39953 => "0000000000101101",39954 => "0000000000101101",
39955 => "0000000000101101",39956 => "0000000000101101",
39957 => "0000000000101101",39958 => "0000000000101101",
39959 => "0000000000101101",39960 => "0000000000101101",
39961 => "0000000000101101",39962 => "0000000000101101",
39963 => "0000000000101101",39964 => "0000000000101101",
39965 => "0000000000101101",39966 => "0000000000101101",
39967 => "0000000000101101",39968 => "0000000000101101",
39969 => "0000000000101101",39970 => "0000000000101101",
39971 => "0000000000101101",39972 => "0000000000101101",
39973 => "0000000000101101",39974 => "0000000000101101",
39975 => "0000000000101101",39976 => "0000000000101101",
39977 => "0000000000101101",39978 => "0000000000101101",
39979 => "0000000000101101",39980 => "0000000000101101",
39981 => "0000000000101101",39982 => "0000000000101101",
39983 => "0000000000101101",39984 => "0000000000101101",
39985 => "0000000000101101",39986 => "0000000000101101",
39987 => "0000000000101101",39988 => "0000000000101101",
39989 => "0000000000101101",39990 => "0000000000101101",
39991 => "0000000000101101",39992 => "0000000000101101",
39993 => "0000000000101101",39994 => "0000000000101101",
39995 => "0000000000101101",39996 => "0000000000101101",
39997 => "0000000000101101",39998 => "0000000000101101",
39999 => "0000000000101101",40000 => "0000000000101101",
40001 => "0000000000101101",40002 => "0000000000101101",
40003 => "0000000000101101",40004 => "0000000000101101",
40005 => "0000000000101101",40006 => "0000000000101101",
40007 => "0000000000101101",40008 => "0000000000101101",
40009 => "0000000000101101",40010 => "0000000000101101",
40011 => "0000000000101101",40012 => "0000000000101101",
40013 => "0000000000101101",40014 => "0000000000101101",
40015 => "0000000000101101",40016 => "0000000000101101",
40017 => "0000000000101101",40018 => "0000000000101101",
40019 => "0000000000101101",40020 => "0000000000101101",
40021 => "0000000000101101",40022 => "0000000000101101",
40023 => "0000000000101101",40024 => "0000000000101101",
40025 => "0000000000101101",40026 => "0000000000101101",
40027 => "0000000000101101",40028 => "0000000000101101",
40029 => "0000000000101101",40030 => "0000000000101101",
40031 => "0000000000101101",40032 => "0000000000101101",
40033 => "0000000000101101",40034 => "0000000000101101",
40035 => "0000000000101100",40036 => "0000000000101100",
40037 => "0000000000101100",40038 => "0000000000101100",
40039 => "0000000000101100",40040 => "0000000000101100",
40041 => "0000000000101100",40042 => "0000000000101100",
40043 => "0000000000101100",40044 => "0000000000101100",
40045 => "0000000000101100",40046 => "0000000000101100",
40047 => "0000000000101100",40048 => "0000000000101100",
40049 => "0000000000101100",40050 => "0000000000101100",
40051 => "0000000000101100",40052 => "0000000000101100",
40053 => "0000000000101100",40054 => "0000000000101100",
40055 => "0000000000101100",40056 => "0000000000101100",
40057 => "0000000000101100",40058 => "0000000000101100",
40059 => "0000000000101100",40060 => "0000000000101100",
40061 => "0000000000101100",40062 => "0000000000101100",
40063 => "0000000000101100",40064 => "0000000000101100",
40065 => "0000000000101100",40066 => "0000000000101100",
40067 => "0000000000101100",40068 => "0000000000101100",
40069 => "0000000000101100",40070 => "0000000000101100",
40071 => "0000000000101100",40072 => "0000000000101100",
40073 => "0000000000101100",40074 => "0000000000101100",
40075 => "0000000000101100",40076 => "0000000000101100",
40077 => "0000000000101100",40078 => "0000000000101100",
40079 => "0000000000101100",40080 => "0000000000101100",
40081 => "0000000000101100",40082 => "0000000000101100",
40083 => "0000000000101100",40084 => "0000000000101100",
40085 => "0000000000101100",40086 => "0000000000101100",
40087 => "0000000000101100",40088 => "0000000000101100",
40089 => "0000000000101100",40090 => "0000000000101100",
40091 => "0000000000101100",40092 => "0000000000101100",
40093 => "0000000000101100",40094 => "0000000000101100",
40095 => "0000000000101100",40096 => "0000000000101100",
40097 => "0000000000101100",40098 => "0000000000101100",
40099 => "0000000000101100",40100 => "0000000000101100",
40101 => "0000000000101100",40102 => "0000000000101100",
40103 => "0000000000101100",40104 => "0000000000101100",
40105 => "0000000000101100",40106 => "0000000000101100",
40107 => "0000000000101100",40108 => "0000000000101100",
40109 => "0000000000101100",40110 => "0000000000101100",
40111 => "0000000000101100",40112 => "0000000000101100",
40113 => "0000000000101100",40114 => "0000000000101100",
40115 => "0000000000101100",40116 => "0000000000101100",
40117 => "0000000000101100",40118 => "0000000000101100",
40119 => "0000000000101100",40120 => "0000000000101100",
40121 => "0000000000101100",40122 => "0000000000101100",
40123 => "0000000000101100",40124 => "0000000000101100",
40125 => "0000000000101100",40126 => "0000000000101100",
40127 => "0000000000101100",40128 => "0000000000101100",
40129 => "0000000000101100",40130 => "0000000000101100",
40131 => "0000000000101100",40132 => "0000000000101100",
40133 => "0000000000101100",40134 => "0000000000101100",
40135 => "0000000000101100",40136 => "0000000000101100",
40137 => "0000000000101100",40138 => "0000000000101100",
40139 => "0000000000101100",40140 => "0000000000101100",
40141 => "0000000000101100",40142 => "0000000000101100",
40143 => "0000000000101100",40144 => "0000000000101100",
40145 => "0000000000101100",40146 => "0000000000101100",
40147 => "0000000000101100",40148 => "0000000000101100",
40149 => "0000000000101100",40150 => "0000000000101100",
40151 => "0000000000101100",40152 => "0000000000101100",
40153 => "0000000000101100",40154 => "0000000000101100",
40155 => "0000000000101100",40156 => "0000000000101100",
40157 => "0000000000101100",40158 => "0000000000101100",
40159 => "0000000000101100",40160 => "0000000000101100",
40161 => "0000000000101100",40162 => "0000000000101100",
40163 => "0000000000101100",40164 => "0000000000101100",
40165 => "0000000000101100",40166 => "0000000000101100",
40167 => "0000000000101100",40168 => "0000000000101100",
40169 => "0000000000101100",40170 => "0000000000101100",
40171 => "0000000000101100",40172 => "0000000000101100",
40173 => "0000000000101100",40174 => "0000000000101100",
40175 => "0000000000101100",40176 => "0000000000101100",
40177 => "0000000000101100",40178 => "0000000000101100",
40179 => "0000000000101100",40180 => "0000000000101100",
40181 => "0000000000101100",40182 => "0000000000101100",
40183 => "0000000000101100",40184 => "0000000000101100",
40185 => "0000000000101100",40186 => "0000000000101100",
40187 => "0000000000101100",40188 => "0000000000101100",
40189 => "0000000000101100",40190 => "0000000000101100",
40191 => "0000000000101100",40192 => "0000000000101100",
40193 => "0000000000101100",40194 => "0000000000101100",
40195 => "0000000000101100",40196 => "0000000000101100",
40197 => "0000000000101100",40198 => "0000000000101100",
40199 => "0000000000101100",40200 => "0000000000101100",
40201 => "0000000000101100",40202 => "0000000000101100",
40203 => "0000000000101100",40204 => "0000000000101100",
40205 => "0000000000101100",40206 => "0000000000101100",
40207 => "0000000000101100",40208 => "0000000000101100",
40209 => "0000000000101100",40210 => "0000000000101100",
40211 => "0000000000101100",40212 => "0000000000101100",
40213 => "0000000000101100",40214 => "0000000000101100",
40215 => "0000000000101100",40216 => "0000000000101100",
40217 => "0000000000101100",40218 => "0000000000101100",
40219 => "0000000000101100",40220 => "0000000000101100",
40221 => "0000000000101100",40222 => "0000000000101100",
40223 => "0000000000101100",40224 => "0000000000101100",
40225 => "0000000000101100",40226 => "0000000000101100",
40227 => "0000000000101100",40228 => "0000000000101100",
40229 => "0000000000101100",40230 => "0000000000101100",
40231 => "0000000000101100",40232 => "0000000000101100",
40233 => "0000000000101100",40234 => "0000000000101100",
40235 => "0000000000101100",40236 => "0000000000101100",
40237 => "0000000000101100",40238 => "0000000000101100",
40239 => "0000000000101100",40240 => "0000000000101100",
40241 => "0000000000101100",40242 => "0000000000101100",
40243 => "0000000000101100",40244 => "0000000000101100",
40245 => "0000000000101100",40246 => "0000000000101100",
40247 => "0000000000101100",40248 => "0000000000101100",
40249 => "0000000000101100",40250 => "0000000000101100",
40251 => "0000000000101100",40252 => "0000000000101100",
40253 => "0000000000101100",40254 => "0000000000101100",
40255 => "0000000000101100",40256 => "0000000000101100",
40257 => "0000000000101100",40258 => "0000000000101100",
40259 => "0000000000101100",40260 => "0000000000101100",
40261 => "0000000000101100",40262 => "0000000000101011",
40263 => "0000000000101011",40264 => "0000000000101011",
40265 => "0000000000101011",40266 => "0000000000101011",
40267 => "0000000000101011",40268 => "0000000000101011",
40269 => "0000000000101011",40270 => "0000000000101011",
40271 => "0000000000101011",40272 => "0000000000101011",
40273 => "0000000000101011",40274 => "0000000000101011",
40275 => "0000000000101011",40276 => "0000000000101011",
40277 => "0000000000101011",40278 => "0000000000101011",
40279 => "0000000000101011",40280 => "0000000000101011",
40281 => "0000000000101011",40282 => "0000000000101011",
40283 => "0000000000101011",40284 => "0000000000101011",
40285 => "0000000000101011",40286 => "0000000000101011",
40287 => "0000000000101011",40288 => "0000000000101011",
40289 => "0000000000101011",40290 => "0000000000101011",
40291 => "0000000000101011",40292 => "0000000000101011",
40293 => "0000000000101011",40294 => "0000000000101011",
40295 => "0000000000101011",40296 => "0000000000101011",
40297 => "0000000000101011",40298 => "0000000000101011",
40299 => "0000000000101011",40300 => "0000000000101011",
40301 => "0000000000101011",40302 => "0000000000101011",
40303 => "0000000000101011",40304 => "0000000000101011",
40305 => "0000000000101011",40306 => "0000000000101011",
40307 => "0000000000101011",40308 => "0000000000101011",
40309 => "0000000000101011",40310 => "0000000000101011",
40311 => "0000000000101011",40312 => "0000000000101011",
40313 => "0000000000101011",40314 => "0000000000101011",
40315 => "0000000000101011",40316 => "0000000000101011",
40317 => "0000000000101011",40318 => "0000000000101011",
40319 => "0000000000101011",40320 => "0000000000101011",
40321 => "0000000000101011",40322 => "0000000000101011",
40323 => "0000000000101011",40324 => "0000000000101011",
40325 => "0000000000101011",40326 => "0000000000101011",
40327 => "0000000000101011",40328 => "0000000000101011",
40329 => "0000000000101011",40330 => "0000000000101011",
40331 => "0000000000101011",40332 => "0000000000101011",
40333 => "0000000000101011",40334 => "0000000000101011",
40335 => "0000000000101011",40336 => "0000000000101011",
40337 => "0000000000101011",40338 => "0000000000101011",
40339 => "0000000000101011",40340 => "0000000000101011",
40341 => "0000000000101011",40342 => "0000000000101011",
40343 => "0000000000101011",40344 => "0000000000101011",
40345 => "0000000000101011",40346 => "0000000000101011",
40347 => "0000000000101011",40348 => "0000000000101011",
40349 => "0000000000101011",40350 => "0000000000101011",
40351 => "0000000000101011",40352 => "0000000000101011",
40353 => "0000000000101011",40354 => "0000000000101011",
40355 => "0000000000101011",40356 => "0000000000101011",
40357 => "0000000000101011",40358 => "0000000000101011",
40359 => "0000000000101011",40360 => "0000000000101011",
40361 => "0000000000101011",40362 => "0000000000101011",
40363 => "0000000000101011",40364 => "0000000000101011",
40365 => "0000000000101011",40366 => "0000000000101011",
40367 => "0000000000101011",40368 => "0000000000101011",
40369 => "0000000000101011",40370 => "0000000000101011",
40371 => "0000000000101011",40372 => "0000000000101011",
40373 => "0000000000101011",40374 => "0000000000101011",
40375 => "0000000000101011",40376 => "0000000000101011",
40377 => "0000000000101011",40378 => "0000000000101011",
40379 => "0000000000101011",40380 => "0000000000101011",
40381 => "0000000000101011",40382 => "0000000000101011",
40383 => "0000000000101011",40384 => "0000000000101011",
40385 => "0000000000101011",40386 => "0000000000101011",
40387 => "0000000000101011",40388 => "0000000000101011",
40389 => "0000000000101011",40390 => "0000000000101011",
40391 => "0000000000101011",40392 => "0000000000101011",
40393 => "0000000000101011",40394 => "0000000000101011",
40395 => "0000000000101011",40396 => "0000000000101011",
40397 => "0000000000101011",40398 => "0000000000101011",
40399 => "0000000000101011",40400 => "0000000000101011",
40401 => "0000000000101011",40402 => "0000000000101011",
40403 => "0000000000101011",40404 => "0000000000101011",
40405 => "0000000000101011",40406 => "0000000000101011",
40407 => "0000000000101011",40408 => "0000000000101011",
40409 => "0000000000101011",40410 => "0000000000101011",
40411 => "0000000000101011",40412 => "0000000000101011",
40413 => "0000000000101011",40414 => "0000000000101011",
40415 => "0000000000101011",40416 => "0000000000101011",
40417 => "0000000000101011",40418 => "0000000000101011",
40419 => "0000000000101011",40420 => "0000000000101011",
40421 => "0000000000101011",40422 => "0000000000101011",
40423 => "0000000000101011",40424 => "0000000000101011",
40425 => "0000000000101011",40426 => "0000000000101011",
40427 => "0000000000101011",40428 => "0000000000101011",
40429 => "0000000000101011",40430 => "0000000000101011",
40431 => "0000000000101011",40432 => "0000000000101011",
40433 => "0000000000101011",40434 => "0000000000101011",
40435 => "0000000000101011",40436 => "0000000000101011",
40437 => "0000000000101011",40438 => "0000000000101011",
40439 => "0000000000101011",40440 => "0000000000101011",
40441 => "0000000000101011",40442 => "0000000000101011",
40443 => "0000000000101011",40444 => "0000000000101011",
40445 => "0000000000101011",40446 => "0000000000101011",
40447 => "0000000000101011",40448 => "0000000000101011",
40449 => "0000000000101011",40450 => "0000000000101011",
40451 => "0000000000101011",40452 => "0000000000101011",
40453 => "0000000000101011",40454 => "0000000000101011",
40455 => "0000000000101011",40456 => "0000000000101011",
40457 => "0000000000101011",40458 => "0000000000101011",
40459 => "0000000000101011",40460 => "0000000000101011",
40461 => "0000000000101011",40462 => "0000000000101011",
40463 => "0000000000101011",40464 => "0000000000101011",
40465 => "0000000000101011",40466 => "0000000000101011",
40467 => "0000000000101011",40468 => "0000000000101011",
40469 => "0000000000101011",40470 => "0000000000101011",
40471 => "0000000000101011",40472 => "0000000000101011",
40473 => "0000000000101011",40474 => "0000000000101011",
40475 => "0000000000101011",40476 => "0000000000101011",
40477 => "0000000000101011",40478 => "0000000000101011",
40479 => "0000000000101011",40480 => "0000000000101011",
40481 => "0000000000101011",40482 => "0000000000101011",
40483 => "0000000000101011",40484 => "0000000000101011",
40485 => "0000000000101011",40486 => "0000000000101011",
40487 => "0000000000101011",40488 => "0000000000101011",
40489 => "0000000000101011",40490 => "0000000000101011",
40491 => "0000000000101011",40492 => "0000000000101011",
40493 => "0000000000101011",40494 => "0000000000101011",
40495 => "0000000000101010",40496 => "0000000000101010",
40497 => "0000000000101010",40498 => "0000000000101010",
40499 => "0000000000101010",40500 => "0000000000101010",
40501 => "0000000000101010",40502 => "0000000000101010",
40503 => "0000000000101010",40504 => "0000000000101010",
40505 => "0000000000101010",40506 => "0000000000101010",
40507 => "0000000000101010",40508 => "0000000000101010",
40509 => "0000000000101010",40510 => "0000000000101010",
40511 => "0000000000101010",40512 => "0000000000101010",
40513 => "0000000000101010",40514 => "0000000000101010",
40515 => "0000000000101010",40516 => "0000000000101010",
40517 => "0000000000101010",40518 => "0000000000101010",
40519 => "0000000000101010",40520 => "0000000000101010",
40521 => "0000000000101010",40522 => "0000000000101010",
40523 => "0000000000101010",40524 => "0000000000101010",
40525 => "0000000000101010",40526 => "0000000000101010",
40527 => "0000000000101010",40528 => "0000000000101010",
40529 => "0000000000101010",40530 => "0000000000101010",
40531 => "0000000000101010",40532 => "0000000000101010",
40533 => "0000000000101010",40534 => "0000000000101010",
40535 => "0000000000101010",40536 => "0000000000101010",
40537 => "0000000000101010",40538 => "0000000000101010",
40539 => "0000000000101010",40540 => "0000000000101010",
40541 => "0000000000101010",40542 => "0000000000101010",
40543 => "0000000000101010",40544 => "0000000000101010",
40545 => "0000000000101010",40546 => "0000000000101010",
40547 => "0000000000101010",40548 => "0000000000101010",
40549 => "0000000000101010",40550 => "0000000000101010",
40551 => "0000000000101010",40552 => "0000000000101010",
40553 => "0000000000101010",40554 => "0000000000101010",
40555 => "0000000000101010",40556 => "0000000000101010",
40557 => "0000000000101010",40558 => "0000000000101010",
40559 => "0000000000101010",40560 => "0000000000101010",
40561 => "0000000000101010",40562 => "0000000000101010",
40563 => "0000000000101010",40564 => "0000000000101010",
40565 => "0000000000101010",40566 => "0000000000101010",
40567 => "0000000000101010",40568 => "0000000000101010",
40569 => "0000000000101010",40570 => "0000000000101010",
40571 => "0000000000101010",40572 => "0000000000101010",
40573 => "0000000000101010",40574 => "0000000000101010",
40575 => "0000000000101010",40576 => "0000000000101010",
40577 => "0000000000101010",40578 => "0000000000101010",
40579 => "0000000000101010",40580 => "0000000000101010",
40581 => "0000000000101010",40582 => "0000000000101010",
40583 => "0000000000101010",40584 => "0000000000101010",
40585 => "0000000000101010",40586 => "0000000000101010",
40587 => "0000000000101010",40588 => "0000000000101010",
40589 => "0000000000101010",40590 => "0000000000101010",
40591 => "0000000000101010",40592 => "0000000000101010",
40593 => "0000000000101010",40594 => "0000000000101010",
40595 => "0000000000101010",40596 => "0000000000101010",
40597 => "0000000000101010",40598 => "0000000000101010",
40599 => "0000000000101010",40600 => "0000000000101010",
40601 => "0000000000101010",40602 => "0000000000101010",
40603 => "0000000000101010",40604 => "0000000000101010",
40605 => "0000000000101010",40606 => "0000000000101010",
40607 => "0000000000101010",40608 => "0000000000101010",
40609 => "0000000000101010",40610 => "0000000000101010",
40611 => "0000000000101010",40612 => "0000000000101010",
40613 => "0000000000101010",40614 => "0000000000101010",
40615 => "0000000000101010",40616 => "0000000000101010",
40617 => "0000000000101010",40618 => "0000000000101010",
40619 => "0000000000101010",40620 => "0000000000101010",
40621 => "0000000000101010",40622 => "0000000000101010",
40623 => "0000000000101010",40624 => "0000000000101010",
40625 => "0000000000101010",40626 => "0000000000101010",
40627 => "0000000000101010",40628 => "0000000000101010",
40629 => "0000000000101010",40630 => "0000000000101010",
40631 => "0000000000101010",40632 => "0000000000101010",
40633 => "0000000000101010",40634 => "0000000000101010",
40635 => "0000000000101010",40636 => "0000000000101010",
40637 => "0000000000101010",40638 => "0000000000101010",
40639 => "0000000000101010",40640 => "0000000000101010",
40641 => "0000000000101010",40642 => "0000000000101010",
40643 => "0000000000101010",40644 => "0000000000101010",
40645 => "0000000000101010",40646 => "0000000000101010",
40647 => "0000000000101010",40648 => "0000000000101010",
40649 => "0000000000101010",40650 => "0000000000101010",
40651 => "0000000000101010",40652 => "0000000000101010",
40653 => "0000000000101010",40654 => "0000000000101010",
40655 => "0000000000101010",40656 => "0000000000101010",
40657 => "0000000000101010",40658 => "0000000000101010",
40659 => "0000000000101010",40660 => "0000000000101010",
40661 => "0000000000101010",40662 => "0000000000101010",
40663 => "0000000000101010",40664 => "0000000000101010",
40665 => "0000000000101010",40666 => "0000000000101010",
40667 => "0000000000101010",40668 => "0000000000101010",
40669 => "0000000000101010",40670 => "0000000000101010",
40671 => "0000000000101010",40672 => "0000000000101010",
40673 => "0000000000101010",40674 => "0000000000101010",
40675 => "0000000000101010",40676 => "0000000000101010",
40677 => "0000000000101010",40678 => "0000000000101010",
40679 => "0000000000101010",40680 => "0000000000101010",
40681 => "0000000000101010",40682 => "0000000000101010",
40683 => "0000000000101010",40684 => "0000000000101010",
40685 => "0000000000101010",40686 => "0000000000101010",
40687 => "0000000000101010",40688 => "0000000000101010",
40689 => "0000000000101010",40690 => "0000000000101010",
40691 => "0000000000101010",40692 => "0000000000101010",
40693 => "0000000000101010",40694 => "0000000000101010",
40695 => "0000000000101010",40696 => "0000000000101010",
40697 => "0000000000101010",40698 => "0000000000101010",
40699 => "0000000000101010",40700 => "0000000000101010",
40701 => "0000000000101010",40702 => "0000000000101010",
40703 => "0000000000101010",40704 => "0000000000101010",
40705 => "0000000000101010",40706 => "0000000000101010",
40707 => "0000000000101010",40708 => "0000000000101010",
40709 => "0000000000101010",40710 => "0000000000101010",
40711 => "0000000000101010",40712 => "0000000000101010",
40713 => "0000000000101010",40714 => "0000000000101010",
40715 => "0000000000101010",40716 => "0000000000101010",
40717 => "0000000000101010",40718 => "0000000000101010",
40719 => "0000000000101010",40720 => "0000000000101010",
40721 => "0000000000101010",40722 => "0000000000101010",
40723 => "0000000000101010",40724 => "0000000000101010",
40725 => "0000000000101010",40726 => "0000000000101010",
40727 => "0000000000101010",40728 => "0000000000101010",
40729 => "0000000000101010",40730 => "0000000000101010",
40731 => "0000000000101010",40732 => "0000000000101010",
40733 => "0000000000101001",40734 => "0000000000101001",
40735 => "0000000000101001",40736 => "0000000000101001",
40737 => "0000000000101001",40738 => "0000000000101001",
40739 => "0000000000101001",40740 => "0000000000101001",
40741 => "0000000000101001",40742 => "0000000000101001",
40743 => "0000000000101001",40744 => "0000000000101001",
40745 => "0000000000101001",40746 => "0000000000101001",
40747 => "0000000000101001",40748 => "0000000000101001",
40749 => "0000000000101001",40750 => "0000000000101001",
40751 => "0000000000101001",40752 => "0000000000101001",
40753 => "0000000000101001",40754 => "0000000000101001",
40755 => "0000000000101001",40756 => "0000000000101001",
40757 => "0000000000101001",40758 => "0000000000101001",
40759 => "0000000000101001",40760 => "0000000000101001",
40761 => "0000000000101001",40762 => "0000000000101001",
40763 => "0000000000101001",40764 => "0000000000101001",
40765 => "0000000000101001",40766 => "0000000000101001",
40767 => "0000000000101001",40768 => "0000000000101001",
40769 => "0000000000101001",40770 => "0000000000101001",
40771 => "0000000000101001",40772 => "0000000000101001",
40773 => "0000000000101001",40774 => "0000000000101001",
40775 => "0000000000101001",40776 => "0000000000101001",
40777 => "0000000000101001",40778 => "0000000000101001",
40779 => "0000000000101001",40780 => "0000000000101001",
40781 => "0000000000101001",40782 => "0000000000101001",
40783 => "0000000000101001",40784 => "0000000000101001",
40785 => "0000000000101001",40786 => "0000000000101001",
40787 => "0000000000101001",40788 => "0000000000101001",
40789 => "0000000000101001",40790 => "0000000000101001",
40791 => "0000000000101001",40792 => "0000000000101001",
40793 => "0000000000101001",40794 => "0000000000101001",
40795 => "0000000000101001",40796 => "0000000000101001",
40797 => "0000000000101001",40798 => "0000000000101001",
40799 => "0000000000101001",40800 => "0000000000101001",
40801 => "0000000000101001",40802 => "0000000000101001",
40803 => "0000000000101001",40804 => "0000000000101001",
40805 => "0000000000101001",40806 => "0000000000101001",
40807 => "0000000000101001",40808 => "0000000000101001",
40809 => "0000000000101001",40810 => "0000000000101001",
40811 => "0000000000101001",40812 => "0000000000101001",
40813 => "0000000000101001",40814 => "0000000000101001",
40815 => "0000000000101001",40816 => "0000000000101001",
40817 => "0000000000101001",40818 => "0000000000101001",
40819 => "0000000000101001",40820 => "0000000000101001",
40821 => "0000000000101001",40822 => "0000000000101001",
40823 => "0000000000101001",40824 => "0000000000101001",
40825 => "0000000000101001",40826 => "0000000000101001",
40827 => "0000000000101001",40828 => "0000000000101001",
40829 => "0000000000101001",40830 => "0000000000101001",
40831 => "0000000000101001",40832 => "0000000000101001",
40833 => "0000000000101001",40834 => "0000000000101001",
40835 => "0000000000101001",40836 => "0000000000101001",
40837 => "0000000000101001",40838 => "0000000000101001",
40839 => "0000000000101001",40840 => "0000000000101001",
40841 => "0000000000101001",40842 => "0000000000101001",
40843 => "0000000000101001",40844 => "0000000000101001",
40845 => "0000000000101001",40846 => "0000000000101001",
40847 => "0000000000101001",40848 => "0000000000101001",
40849 => "0000000000101001",40850 => "0000000000101001",
40851 => "0000000000101001",40852 => "0000000000101001",
40853 => "0000000000101001",40854 => "0000000000101001",
40855 => "0000000000101001",40856 => "0000000000101001",
40857 => "0000000000101001",40858 => "0000000000101001",
40859 => "0000000000101001",40860 => "0000000000101001",
40861 => "0000000000101001",40862 => "0000000000101001",
40863 => "0000000000101001",40864 => "0000000000101001",
40865 => "0000000000101001",40866 => "0000000000101001",
40867 => "0000000000101001",40868 => "0000000000101001",
40869 => "0000000000101001",40870 => "0000000000101001",
40871 => "0000000000101001",40872 => "0000000000101001",
40873 => "0000000000101001",40874 => "0000000000101001",
40875 => "0000000000101001",40876 => "0000000000101001",
40877 => "0000000000101001",40878 => "0000000000101001",
40879 => "0000000000101001",40880 => "0000000000101001",
40881 => "0000000000101001",40882 => "0000000000101001",
40883 => "0000000000101001",40884 => "0000000000101001",
40885 => "0000000000101001",40886 => "0000000000101001",
40887 => "0000000000101001",40888 => "0000000000101001",
40889 => "0000000000101001",40890 => "0000000000101001",
40891 => "0000000000101001",40892 => "0000000000101001",
40893 => "0000000000101001",40894 => "0000000000101001",
40895 => "0000000000101001",40896 => "0000000000101001",
40897 => "0000000000101001",40898 => "0000000000101001",
40899 => "0000000000101001",40900 => "0000000000101001",
40901 => "0000000000101001",40902 => "0000000000101001",
40903 => "0000000000101001",40904 => "0000000000101001",
40905 => "0000000000101001",40906 => "0000000000101001",
40907 => "0000000000101001",40908 => "0000000000101001",
40909 => "0000000000101001",40910 => "0000000000101001",
40911 => "0000000000101001",40912 => "0000000000101001",
40913 => "0000000000101001",40914 => "0000000000101001",
40915 => "0000000000101001",40916 => "0000000000101001",
40917 => "0000000000101001",40918 => "0000000000101001",
40919 => "0000000000101001",40920 => "0000000000101001",
40921 => "0000000000101001",40922 => "0000000000101001",
40923 => "0000000000101001",40924 => "0000000000101001",
40925 => "0000000000101001",40926 => "0000000000101001",
40927 => "0000000000101001",40928 => "0000000000101001",
40929 => "0000000000101001",40930 => "0000000000101001",
40931 => "0000000000101001",40932 => "0000000000101001",
40933 => "0000000000101001",40934 => "0000000000101001",
40935 => "0000000000101001",40936 => "0000000000101001",
40937 => "0000000000101001",40938 => "0000000000101001",
40939 => "0000000000101001",40940 => "0000000000101001",
40941 => "0000000000101001",40942 => "0000000000101001",
40943 => "0000000000101001",40944 => "0000000000101001",
40945 => "0000000000101001",40946 => "0000000000101001",
40947 => "0000000000101001",40948 => "0000000000101001",
40949 => "0000000000101001",40950 => "0000000000101001",
40951 => "0000000000101001",40952 => "0000000000101001",
40953 => "0000000000101001",40954 => "0000000000101001",
40955 => "0000000000101001",40956 => "0000000000101001",
40957 => "0000000000101001",40958 => "0000000000101001",
40959 => "0000000000101001",40960 => "0000000000010010",
40961 => "0000000000010001",40962 => "0000000000001111",
40963 => "0000000000001110",40964 => "0000000000001100",
40965 => "0000000000001011",40966 => "0000000000000001",
40967 => "0000000000001001",40968 => "0000000000001000",
40969 => "0000000000000111",40970 => "0000000000010001",
40971 => "0000000000010000",40972 => "0000000000010000",
40973 => "0000000000010000",40974 => "0000000000010000",
40975 => "0000000000010000",40976 => "0000000000010000",
40977 => "0000000000001111",40978 => "0000000000001111",
40979 => "0000000000001111",40980 => "0000000000001111",
40981 => "0000000000001111",40982 => "0000000000001111",
40983 => "0000000000001111",40984 => "0000000000001110",
40985 => "0000000000001110",40986 => "0000000000001110",
40987 => "0000000000001110",40988 => "0000000000001110",
40989 => "0000000000001110",40990 => "0000000000001110",
40991 => "0000000000001101",40992 => "0000000000001101",
40993 => "0000000000001101",40994 => "0000000000001101",
40995 => "0000000000001101",40996 => "0000000000001101",
40997 => "0000000000001101",40998 => "0000000000001101",
40999 => "0000000000001100",41000 => "0000000000001100",
41001 => "0000000000001100",41002 => "0000000000001100",
41003 => "0000000000001100",41004 => "0000000000001100",
41005 => "0000000000001100",41006 => "0000000000001100",
41007 => "0000000000001011",41008 => "0000000000001011",
41009 => "0000000000001011",41010 => "0000000000001011",
41011 => "0000000000001011",41012 => "0000000000001011",
41013 => "0000000000001011",41014 => "0000000000001011",
41015 => "0000000000001011",41016 => "0000000000000001",
41017 => "0000000000000001",41018 => "0000000000000001",
41019 => "0000000000000001",41020 => "0000000000000001",
41021 => "0000000000000001",41022 => "0000000000000001",
41023 => "0000000000000001",41024 => "0000000000000001",
41025 => "0000000000000001",41026 => "0000000000001001",
41027 => "0000000000001001",41028 => "0000000000001001",
41029 => "0000000000001001",41030 => "0000000000001001",
41031 => "0000000000001001",41032 => "0000000000001001",
41033 => "0000000000001001",41034 => "0000000000001001",
41035 => "0000000000001001",41036 => "0000000000001001",
41037 => "0000000000001000",41038 => "0000000000001000",
41039 => "0000000000001000",41040 => "0000000000001000",
41041 => "0000000000001000",41042 => "0000000000001000",
41043 => "0000000000001000",41044 => "0000000000001000",
41045 => "0000000000001000",41046 => "0000000000001000",
41047 => "0000000000001000",41048 => "0000000000001000",
41049 => "0000000000001000",41050 => "0000000000000111",
41051 => "0000000000000111",41052 => "0000000000000111",
41053 => "0000000000000111",41054 => "0000000000000111",
41055 => "0000000000000111",41056 => "0000000000000111",
41057 => "0000000000000111",41058 => "0000000000000111",
41059 => "0000000000000111",41060 => "0000000000010001",
41061 => "0000000000010001",41062 => "0000000000010001",
41063 => "0000000000010001",41064 => "0000000000010001",
41065 => "0000000000010000",41066 => "0000000000010000",
41067 => "0000000000010000",41068 => "0000000000010000",
41069 => "0000000000010000",41070 => "0000000000010000",
41071 => "0000000000010000",41072 => "0000000000010000",
41073 => "0000000000010000",41074 => "0000000000010000",
41075 => "0000000000010000",41076 => "0000000000010000",
41077 => "0000000000010000",41078 => "0000000000010000",
41079 => "0000000000010000",41080 => "0000000000010000",
41081 => "0000000000010000",41082 => "0000000000010000",
41083 => "0000000000010000",41084 => "0000000000010000",
41085 => "0000000000010000",41086 => "0000000000010000",
41087 => "0000000000010000",41088 => "0000000000010000",
41089 => "0000000000010000",41090 => "0000000000010000",
41091 => "0000000000010000",41092 => "0000000000010000",
41093 => "0000000000010000",41094 => "0000000000010000",
41095 => "0000000000010000",41096 => "0000000000010000",
41097 => "0000000000010000",41098 => "0000000000010000",
41099 => "0000000000010000",41100 => "0000000000010000",
41101 => "0000000000010000",41102 => "0000000000010000",
41103 => "0000000000010000",41104 => "0000000000010000",
41105 => "0000000000010000",41106 => "0000000000010000",
41107 => "0000000000010000",41108 => "0000000000010000",
41109 => "0000000000010000",41110 => "0000000000010000",
41111 => "0000000000010000",41112 => "0000000000010000",
41113 => "0000000000010000",41114 => "0000000000010000",
41115 => "0000000000010000",41116 => "0000000000010000",
41117 => "0000000000010000",41118 => "0000000000010000",
41119 => "0000000000010000",41120 => "0000000000010000",
41121 => "0000000000010000",41122 => "0000000000010000",
41123 => "0000000000010000",41124 => "0000000000010000",
41125 => "0000000000010000",41126 => "0000000000010000",
41127 => "0000000000001111",41128 => "0000000000001111",
41129 => "0000000000001111",41130 => "0000000000001111",
41131 => "0000000000001111",41132 => "0000000000001111",
41133 => "0000000000001111",41134 => "0000000000001111",
41135 => "0000000000001111",41136 => "0000000000001111",
41137 => "0000000000001111",41138 => "0000000000001111",
41139 => "0000000000001111",41140 => "0000000000001111",
41141 => "0000000000001111",41142 => "0000000000001111",
41143 => "0000000000001111",41144 => "0000000000001111",
41145 => "0000000000001111",41146 => "0000000000001111",
41147 => "0000000000001111",41148 => "0000000000001111",
41149 => "0000000000001111",41150 => "0000000000001111",
41151 => "0000000000001111",41152 => "0000000000001111",
41153 => "0000000000001111",41154 => "0000000000001111",
41155 => "0000000000001111",41156 => "0000000000001111",
41157 => "0000000000001111",41158 => "0000000000001111",
41159 => "0000000000001111",41160 => "0000000000001111",
41161 => "0000000000001111",41162 => "0000000000001111",
41163 => "0000000000001111",41164 => "0000000000001111",
41165 => "0000000000001111",41166 => "0000000000001111",
41167 => "0000000000001111",41168 => "0000000000001111",
41169 => "0000000000001111",41170 => "0000000000001111",
41171 => "0000000000001111",41172 => "0000000000001111",
41173 => "0000000000001111",41174 => "0000000000001111",
41175 => "0000000000001111",41176 => "0000000000001111",
41177 => "0000000000001111",41178 => "0000000000001111",
41179 => "0000000000001111",41180 => "0000000000001111",
41181 => "0000000000001111",41182 => "0000000000001111",
41183 => "0000000000001111",41184 => "0000000000001111",
41185 => "0000000000001111",41186 => "0000000000001111",
41187 => "0000000000001111",41188 => "0000000000001111",
41189 => "0000000000001111",41190 => "0000000000001111",
41191 => "0000000000001111",41192 => "0000000000001111",
41193 => "0000000000001111",41194 => "0000000000001110",
41195 => "0000000000001110",41196 => "0000000000001110",
41197 => "0000000000001110",41198 => "0000000000001110",
41199 => "0000000000001110",41200 => "0000000000001110",
41201 => "0000000000001110",41202 => "0000000000001110",
41203 => "0000000000001110",41204 => "0000000000001110",
41205 => "0000000000001110",41206 => "0000000000001110",
41207 => "0000000000001110",41208 => "0000000000001110",
41209 => "0000000000001110",41210 => "0000000000001110",
41211 => "0000000000001110",41212 => "0000000000001110",
41213 => "0000000000001110",41214 => "0000000000001110",
41215 => "0000000000001110",41216 => "0000000000001110",
41217 => "0000000000001110",41218 => "0000000000001110",
41219 => "0000000000001110",41220 => "0000000000001110",
41221 => "0000000000001110",41222 => "0000000000001110",
41223 => "0000000000001110",41224 => "0000000000001110",
41225 => "0000000000001110",41226 => "0000000000001110",
41227 => "0000000000001110",41228 => "0000000000001110",
41229 => "0000000000001110",41230 => "0000000000001110",
41231 => "0000000000001110",41232 => "0000000000001110",
41233 => "0000000000001110",41234 => "0000000000001110",
41235 => "0000000000001110",41236 => "0000000000001110",
41237 => "0000000000001110",41238 => "0000000000001110",
41239 => "0000000000001110",41240 => "0000000000001110",
41241 => "0000000000001110",41242 => "0000000000001110",
41243 => "0000000000001110",41244 => "0000000000001110",
41245 => "0000000000001110",41246 => "0000000000001110",
41247 => "0000000000001110",41248 => "0000000000001110",
41249 => "0000000000001110",41250 => "0000000000001110",
41251 => "0000000000001110",41252 => "0000000000001110",
41253 => "0000000000001110",41254 => "0000000000001110",
41255 => "0000000000001110",41256 => "0000000000001110",
41257 => "0000000000001110",41258 => "0000000000001110",
41259 => "0000000000001110",41260 => "0000000000001110",
41261 => "0000000000001110",41262 => "0000000000001110",
41263 => "0000000000001110",41264 => "0000000000001110",
41265 => "0000000000001110",41266 => "0000000000001101",
41267 => "0000000000001101",41268 => "0000000000001101",
41269 => "0000000000001101",41270 => "0000000000001101",
41271 => "0000000000001101",41272 => "0000000000001101",
41273 => "0000000000001101",41274 => "0000000000001101",
41275 => "0000000000001101",41276 => "0000000000001101",
41277 => "0000000000001101",41278 => "0000000000001101",
41279 => "0000000000001101",41280 => "0000000000001101",
41281 => "0000000000001101",41282 => "0000000000001101",
41283 => "0000000000001101",41284 => "0000000000001101",
41285 => "0000000000001101",41286 => "0000000000001101",
41287 => "0000000000001101",41288 => "0000000000001101",
41289 => "0000000000001101",41290 => "0000000000001101",
41291 => "0000000000001101",41292 => "0000000000001101",
41293 => "0000000000001101",41294 => "0000000000001101",
41295 => "0000000000001101",41296 => "0000000000001101",
41297 => "0000000000001101",41298 => "0000000000001101",
41299 => "0000000000001101",41300 => "0000000000001101",
41301 => "0000000000001101",41302 => "0000000000001101",
41303 => "0000000000001101",41304 => "0000000000001101",
41305 => "0000000000001101",41306 => "0000000000001101",
41307 => "0000000000001101",41308 => "0000000000001101",
41309 => "0000000000001101",41310 => "0000000000001101",
41311 => "0000000000001101",41312 => "0000000000001101",
41313 => "0000000000001101",41314 => "0000000000001101",
41315 => "0000000000001101",41316 => "0000000000001101",
41317 => "0000000000001101",41318 => "0000000000001101",
41319 => "0000000000001101",41320 => "0000000000001101",
41321 => "0000000000001101",41322 => "0000000000001101",
41323 => "0000000000001101",41324 => "0000000000001101",
41325 => "0000000000001101",41326 => "0000000000001101",
41327 => "0000000000001101",41328 => "0000000000001101",
41329 => "0000000000001101",41330 => "0000000000001101",
41331 => "0000000000001101",41332 => "0000000000001101",
41333 => "0000000000001101",41334 => "0000000000001101",
41335 => "0000000000001101",41336 => "0000000000001101",
41337 => "0000000000001101",41338 => "0000000000001101",
41339 => "0000000000001101",41340 => "0000000000001101",
41341 => "0000000000001101",41342 => "0000000000001101",
41343 => "0000000000001100",41344 => "0000000000001100",
41345 => "0000000000001100",41346 => "0000000000001100",
41347 => "0000000000001100",41348 => "0000000000001100",
41349 => "0000000000001100",41350 => "0000000000001100",
41351 => "0000000000001100",41352 => "0000000000001100",
41353 => "0000000000001100",41354 => "0000000000001100",
41355 => "0000000000001100",41356 => "0000000000001100",
41357 => "0000000000001100",41358 => "0000000000001100",
41359 => "0000000000001100",41360 => "0000000000001100",
41361 => "0000000000001100",41362 => "0000000000001100",
41363 => "0000000000001100",41364 => "0000000000001100",
41365 => "0000000000001100",41366 => "0000000000001100",
41367 => "0000000000001100",41368 => "0000000000001100",
41369 => "0000000000001100",41370 => "0000000000001100",
41371 => "0000000000001100",41372 => "0000000000001100",
41373 => "0000000000001100",41374 => "0000000000001100",
41375 => "0000000000001100",41376 => "0000000000001100",
41377 => "0000000000001100",41378 => "0000000000001100",
41379 => "0000000000001100",41380 => "0000000000001100",
41381 => "0000000000001100",41382 => "0000000000001100",
41383 => "0000000000001100",41384 => "0000000000001100",
41385 => "0000000000001100",41386 => "0000000000001100",
41387 => "0000000000001100",41388 => "0000000000001100",
41389 => "0000000000001100",41390 => "0000000000001100",
41391 => "0000000000001100",41392 => "0000000000001100",
41393 => "0000000000001100",41394 => "0000000000001100",
41395 => "0000000000001100",41396 => "0000000000001100",
41397 => "0000000000001100",41398 => "0000000000001100",
41399 => "0000000000001100",41400 => "0000000000001100",
41401 => "0000000000001100",41402 => "0000000000001100",
41403 => "0000000000001100",41404 => "0000000000001100",
41405 => "0000000000001100",41406 => "0000000000001100",
41407 => "0000000000001100",41408 => "0000000000001100",
41409 => "0000000000001100",41410 => "0000000000001100",
41411 => "0000000000001100",41412 => "0000000000001100",
41413 => "0000000000001100",41414 => "0000000000001100",
41415 => "0000000000001100",41416 => "0000000000001100",
41417 => "0000000000001100",41418 => "0000000000001100",
41419 => "0000000000001100",41420 => "0000000000001100",
41421 => "0000000000001100",41422 => "0000000000001100",
41423 => "0000000000001100",41424 => "0000000000001100",
41425 => "0000000000001100",41426 => "0000000000001011",
41427 => "0000000000001011",41428 => "0000000000001011",
41429 => "0000000000001011",41430 => "0000000000001011",
41431 => "0000000000001011",41432 => "0000000000001011",
41433 => "0000000000001011",41434 => "0000000000001011",
41435 => "0000000000001011",41436 => "0000000000001011",
41437 => "0000000000001011",41438 => "0000000000001011",
41439 => "0000000000001011",41440 => "0000000000001011",
41441 => "0000000000001011",41442 => "0000000000001011",
41443 => "0000000000001011",41444 => "0000000000001011",
41445 => "0000000000001011",41446 => "0000000000001011",
41447 => "0000000000001011",41448 => "0000000000001011",
41449 => "0000000000001011",41450 => "0000000000001011",
41451 => "0000000000001011",41452 => "0000000000001011",
41453 => "0000000000001011",41454 => "0000000000001011",
41455 => "0000000000001011",41456 => "0000000000001011",
41457 => "0000000000001011",41458 => "0000000000001011",
41459 => "0000000000001011",41460 => "0000000000001011",
41461 => "0000000000001011",41462 => "0000000000001011",
41463 => "0000000000001011",41464 => "0000000000001011",
41465 => "0000000000001011",41466 => "0000000000001011",
41467 => "0000000000001011",41468 => "0000000000001011",
41469 => "0000000000001011",41470 => "0000000000001011",
41471 => "0000000000001011",41472 => "0000000000001011",
41473 => "0000000000001011",41474 => "0000000000001011",
41475 => "0000000000001011",41476 => "0000000000001011",
41477 => "0000000000001011",41478 => "0000000000001011",
41479 => "0000000000001011",41480 => "0000000000001011",
41481 => "0000000000001011",41482 => "0000000000001011",
41483 => "0000000000001011",41484 => "0000000000001011",
41485 => "0000000000001011",41486 => "0000000000001011",
41487 => "0000000000001011",41488 => "0000000000001011",
41489 => "0000000000001011",41490 => "0000000000001011",
41491 => "0000000000001011",41492 => "0000000000001011",
41493 => "0000000000001011",41494 => "0000000000001011",
41495 => "0000000000001011",41496 => "0000000000001011",
41497 => "0000000000001011",41498 => "0000000000001011",
41499 => "0000000000001011",41500 => "0000000000001011",
41501 => "0000000000001011",41502 => "0000000000001011",
41503 => "0000000000001011",41504 => "0000000000001011",
41505 => "0000000000001011",41506 => "0000000000001011",
41507 => "0000000000001011",41508 => "0000000000001011",
41509 => "0000000000001011",41510 => "0000000000001011",
41511 => "0000000000001011",41512 => "0000000000001011",
41513 => "0000000000001011",41514 => "0000000000001011",
41515 => "0000000000001011",41516 => "0000000000001011",
41517 => "0000000000000001",41518 => "0000000000000001",
41519 => "0000000000000001",41520 => "0000000000000001",
41521 => "0000000000000001",41522 => "0000000000000001",
41523 => "0000000000000001",41524 => "0000000000000001",
41525 => "0000000000000001",41526 => "0000000000000001",
41527 => "0000000000000001",41528 => "0000000000000001",
41529 => "0000000000000001",41530 => "0000000000000001",
41531 => "0000000000000001",41532 => "0000000000000001",
41533 => "0000000000000001",41534 => "0000000000000001",
41535 => "0000000000000001",41536 => "0000000000000001",
41537 => "0000000000000001",41538 => "0000000000000001",
41539 => "0000000000000001",41540 => "0000000000000001",
41541 => "0000000000000001",41542 => "0000000000000001",
41543 => "0000000000000001",41544 => "0000000000000001",
41545 => "0000000000000001",41546 => "0000000000000001",
41547 => "0000000000000001",41548 => "0000000000000001",
41549 => "0000000000000001",41550 => "0000000000000001",
41551 => "0000000000000001",41552 => "0000000000000001",
41553 => "0000000000000001",41554 => "0000000000000001",
41555 => "0000000000000001",41556 => "0000000000000001",
41557 => "0000000000000001",41558 => "0000000000000001",
41559 => "0000000000000001",41560 => "0000000000000001",
41561 => "0000000000000001",41562 => "0000000000000001",
41563 => "0000000000000001",41564 => "0000000000000001",
41565 => "0000000000000001",41566 => "0000000000000001",
41567 => "0000000000000001",41568 => "0000000000000001",
41569 => "0000000000000001",41570 => "0000000000000001",
41571 => "0000000000000001",41572 => "0000000000000001",
41573 => "0000000000000001",41574 => "0000000000000001",
41575 => "0000000000000001",41576 => "0000000000000001",
41577 => "0000000000000001",41578 => "0000000000000001",
41579 => "0000000000000001",41580 => "0000000000000001",
41581 => "0000000000000001",41582 => "0000000000000001",
41583 => "0000000000000001",41584 => "0000000000000001",
41585 => "0000000000000001",41586 => "0000000000000001",
41587 => "0000000000000001",41588 => "0000000000000001",
41589 => "0000000000000001",41590 => "0000000000000001",
41591 => "0000000000000001",41592 => "0000000000000001",
41593 => "0000000000000001",41594 => "0000000000000001",
41595 => "0000000000000001",41596 => "0000000000000001",
41597 => "0000000000000001",41598 => "0000000000000001",
41599 => "0000000000000001",41600 => "0000000000000001",
41601 => "0000000000000001",41602 => "0000000000000001",
41603 => "0000000000000001",41604 => "0000000000000001",
41605 => "0000000000000001",41606 => "0000000000000001",
41607 => "0000000000000001",41608 => "0000000000000001",
41609 => "0000000000000001",41610 => "0000000000000001",
41611 => "0000000000000001",41612 => "0000000000000001",
41613 => "0000000000000001",41614 => "0000000000000001",
41615 => "0000000000000001",41616 => "0000000000000001",
41617 => "0000000000001001",41618 => "0000000000001001",
41619 => "0000000000001001",41620 => "0000000000001001",
41621 => "0000000000001001",41622 => "0000000000001001",
41623 => "0000000000001001",41624 => "0000000000001001",
41625 => "0000000000001001",41626 => "0000000000001001",
41627 => "0000000000001001",41628 => "0000000000001001",
41629 => "0000000000001001",41630 => "0000000000001001",
41631 => "0000000000001001",41632 => "0000000000001001",
41633 => "0000000000001001",41634 => "0000000000001001",
41635 => "0000000000001001",41636 => "0000000000001001",
41637 => "0000000000001001",41638 => "0000000000001001",
41639 => "0000000000001001",41640 => "0000000000001001",
41641 => "0000000000001001",41642 => "0000000000001001",
41643 => "0000000000001001",41644 => "0000000000001001",
41645 => "0000000000001001",41646 => "0000000000001001",
41647 => "0000000000001001",41648 => "0000000000001001",
41649 => "0000000000001001",41650 => "0000000000001001",
41651 => "0000000000001001",41652 => "0000000000001001",
41653 => "0000000000001001",41654 => "0000000000001001",
41655 => "0000000000001001",41656 => "0000000000001001",
41657 => "0000000000001001",41658 => "0000000000001001",
41659 => "0000000000001001",41660 => "0000000000001001",
41661 => "0000000000001001",41662 => "0000000000001001",
41663 => "0000000000001001",41664 => "0000000000001001",
41665 => "0000000000001001",41666 => "0000000000001001",
41667 => "0000000000001001",41668 => "0000000000001001",
41669 => "0000000000001001",41670 => "0000000000001001",
41671 => "0000000000001001",41672 => "0000000000001001",
41673 => "0000000000001001",41674 => "0000000000001001",
41675 => "0000000000001001",41676 => "0000000000001001",
41677 => "0000000000001001",41678 => "0000000000001001",
41679 => "0000000000001001",41680 => "0000000000001001",
41681 => "0000000000001001",41682 => "0000000000001001",
41683 => "0000000000001001",41684 => "0000000000001001",
41685 => "0000000000001001",41686 => "0000000000001001",
41687 => "0000000000001001",41688 => "0000000000001001",
41689 => "0000000000001001",41690 => "0000000000001001",
41691 => "0000000000001001",41692 => "0000000000001001",
41693 => "0000000000001001",41694 => "0000000000001001",
41695 => "0000000000001001",41696 => "0000000000001001",
41697 => "0000000000001001",41698 => "0000000000001001",
41699 => "0000000000001001",41700 => "0000000000001001",
41701 => "0000000000001001",41702 => "0000000000001001",
41703 => "0000000000001001",41704 => "0000000000001001",
41705 => "0000000000001001",41706 => "0000000000001001",
41707 => "0000000000001001",41708 => "0000000000001001",
41709 => "0000000000001001",41710 => "0000000000001001",
41711 => "0000000000001001",41712 => "0000000000001001",
41713 => "0000000000001001",41714 => "0000000000001001",
41715 => "0000000000001001",41716 => "0000000000001001",
41717 => "0000000000001001",41718 => "0000000000001001",
41719 => "0000000000001001",41720 => "0000000000001001",
41721 => "0000000000001001",41722 => "0000000000001001",
41723 => "0000000000001001",41724 => "0000000000001001",
41725 => "0000000000001001",41726 => "0000000000001001",
41727 => "0000000000001001",41728 => "0000000000001000",
41729 => "0000000000001000",41730 => "0000000000001000",
41731 => "0000000000001000",41732 => "0000000000001000",
41733 => "0000000000001000",41734 => "0000000000001000",
41735 => "0000000000001000",41736 => "0000000000001000",
41737 => "0000000000001000",41738 => "0000000000001000",
41739 => "0000000000001000",41740 => "0000000000001000",
41741 => "0000000000001000",41742 => "0000000000001000",
41743 => "0000000000001000",41744 => "0000000000001000",
41745 => "0000000000001000",41746 => "0000000000001000",
41747 => "0000000000001000",41748 => "0000000000001000",
41749 => "0000000000001000",41750 => "0000000000001000",
41751 => "0000000000001000",41752 => "0000000000001000",
41753 => "0000000000001000",41754 => "0000000000001000",
41755 => "0000000000001000",41756 => "0000000000001000",
41757 => "0000000000001000",41758 => "0000000000001000",
41759 => "0000000000001000",41760 => "0000000000001000",
41761 => "0000000000001000",41762 => "0000000000001000",
41763 => "0000000000001000",41764 => "0000000000001000",
41765 => "0000000000001000",41766 => "0000000000001000",
41767 => "0000000000001000",41768 => "0000000000001000",
41769 => "0000000000001000",41770 => "0000000000001000",
41771 => "0000000000001000",41772 => "0000000000001000",
41773 => "0000000000001000",41774 => "0000000000001000",
41775 => "0000000000001000",41776 => "0000000000001000",
41777 => "0000000000001000",41778 => "0000000000001000",
41779 => "0000000000001000",41780 => "0000000000001000",
41781 => "0000000000001000",41782 => "0000000000001000",
41783 => "0000000000001000",41784 => "0000000000001000",
41785 => "0000000000001000",41786 => "0000000000001000",
41787 => "0000000000001000",41788 => "0000000000001000",
41789 => "0000000000001000",41790 => "0000000000001000",
41791 => "0000000000001000",41792 => "0000000000001000",
41793 => "0000000000001000",41794 => "0000000000001000",
41795 => "0000000000001000",41796 => "0000000000001000",
41797 => "0000000000001000",41798 => "0000000000001000",
41799 => "0000000000001000",41800 => "0000000000001000",
41801 => "0000000000001000",41802 => "0000000000001000",
41803 => "0000000000001000",41804 => "0000000000001000",
41805 => "0000000000001000",41806 => "0000000000001000",
41807 => "0000000000001000",41808 => "0000000000001000",
41809 => "0000000000001000",41810 => "0000000000001000",
41811 => "0000000000001000",41812 => "0000000000001000",
41813 => "0000000000001000",41814 => "0000000000001000",
41815 => "0000000000001000",41816 => "0000000000001000",
41817 => "0000000000001000",41818 => "0000000000001000",
41819 => "0000000000001000",41820 => "0000000000001000",
41821 => "0000000000001000",41822 => "0000000000001000",
41823 => "0000000000001000",41824 => "0000000000001000",
41825 => "0000000000001000",41826 => "0000000000001000",
41827 => "0000000000001000",41828 => "0000000000001000",
41829 => "0000000000001000",41830 => "0000000000001000",
41831 => "0000000000001000",41832 => "0000000000001000",
41833 => "0000000000001000",41834 => "0000000000001000",
41835 => "0000000000001000",41836 => "0000000000001000",
41837 => "0000000000001000",41838 => "0000000000001000",
41839 => "0000000000001000",41840 => "0000000000001000",
41841 => "0000000000001000",41842 => "0000000000001000",
41843 => "0000000000001000",41844 => "0000000000001000",
41845 => "0000000000001000",41846 => "0000000000001000",
41847 => "0000000000001000",41848 => "0000000000001000",
41849 => "0000000000001000",41850 => "0000000000001000",
41851 => "0000000000001000",41852 => "0000000000001000",
41853 => "0000000000000111",41854 => "0000000000000111",
41855 => "0000000000000111",41856 => "0000000000000111",
41857 => "0000000000000111",41858 => "0000000000000111",
41859 => "0000000000000111",41860 => "0000000000000111",
41861 => "0000000000000111",41862 => "0000000000000111",
41863 => "0000000000000111",41864 => "0000000000000111",
41865 => "0000000000000111",41866 => "0000000000000111",
41867 => "0000000000000111",41868 => "0000000000000111",
41869 => "0000000000000111",41870 => "0000000000000111",
41871 => "0000000000000111",41872 => "0000000000000111",
41873 => "0000000000000111",41874 => "0000000000000111",
41875 => "0000000000000111",41876 => "0000000000000111",
41877 => "0000000000000111",41878 => "0000000000000111",
41879 => "0000000000000111",41880 => "0000000000000111",
41881 => "0000000000000111",41882 => "0000000000000111",
41883 => "0000000000000111",41884 => "0000000000000111",
41885 => "0000000000000111",41886 => "0000000000000111",
41887 => "0000000000000111",41888 => "0000000000000111",
41889 => "0000000000000111",41890 => "0000000000000111",
41891 => "0000000000000111",41892 => "0000000000000111",
41893 => "0000000000000111",41894 => "0000000000000111",
41895 => "0000000000000111",41896 => "0000000000000111",
41897 => "0000000000000111",41898 => "0000000000000111",
41899 => "0000000000000111",41900 => "0000000000000111",
41901 => "0000000000000111",41902 => "0000000000000111",
41903 => "0000000000000111",41904 => "0000000000000111",
41905 => "0000000000000111",41906 => "0000000000000111",
41907 => "0000000000000111",41908 => "0000000000000111",
41909 => "0000000000000111",41910 => "0000000000000111",
41911 => "0000000000000111",41912 => "0000000000000111",
41913 => "0000000000000111",41914 => "0000000000000111",
41915 => "0000000000000111",41916 => "0000000000000111",
41917 => "0000000000000111",41918 => "0000000000000111",
41919 => "0000000000000111",41920 => "0000000000000111",
41921 => "0000000000000111",41922 => "0000000000000111",
41923 => "0000000000000111",41924 => "0000000000000111",
41925 => "0000000000000111",41926 => "0000000000000111",
41927 => "0000000000000111",41928 => "0000000000000111",
41929 => "0000000000000111",41930 => "0000000000000111",
41931 => "0000000000000111",41932 => "0000000000000111",
41933 => "0000000000000111",41934 => "0000000000000111",
41935 => "0000000000000111",41936 => "0000000000000111",
41937 => "0000000000000111",41938 => "0000000000000111",
41939 => "0000000000000111",41940 => "0000000000000111",
41941 => "0000000000000111",41942 => "0000000000000111",
41943 => "0000000000000111",41944 => "0000000000000111",
41945 => "0000000000000111",41946 => "0000000000000111",
41947 => "0000000000000111",41948 => "0000000000000111",
41949 => "0000000000000111",41950 => "0000000000000111",
41951 => "0000000000000111",41952 => "0000000000000111",
41953 => "0000000000000111",41954 => "0000000000000111",
41955 => "0000000000000111",41956 => "0000000000000111",
41957 => "0000000000000111",41958 => "0000000000000111",
41959 => "0000000000000111",41960 => "0000000000010001",
41961 => "0000000000010001",41962 => "0000000000010001",
41963 => "0000000000010001",41964 => "0000000000010001",
41965 => "0000000000010001",41966 => "0000000000010001",
41967 => "0000000000010001",41968 => "0000000000010001",
41969 => "0000000000010001",41970 => "0000000000010001",
41971 => "0000000000010001",41972 => "0000000000010001",
41973 => "0000000000010001",41974 => "0000000000010001",
41975 => "0000000000010001",41976 => "0000000000010001",
41977 => "0000000000010001",41978 => "0000000000010001",
41979 => "0000000000010001",41980 => "0000000000010001",
41981 => "0000000000010001",41982 => "0000000000010001",
41983 => "0000000000010001",41984 => "0000000000010001",
41985 => "0000000000010001",41986 => "0000000000010001",
41987 => "0000000000010001",41988 => "0000000000010001",
41989 => "0000000000010001",41990 => "0000000000010001",
41991 => "0000000000010001",41992 => "0000000000010001",
41993 => "0000000000010001",41994 => "0000000000010001",
41995 => "0000000000010001",41996 => "0000000000010001",
41997 => "0000000000010001",41998 => "0000000000010001",
41999 => "0000000000010001",42000 => "0000000000010001",
42001 => "0000000000010001",42002 => "0000000000010001",
42003 => "0000000000010001",42004 => "0000000000010000",
42005 => "0000000000010000",42006 => "0000000000010000",
42007 => "0000000000010000",42008 => "0000000000010000",
42009 => "0000000000010000",42010 => "0000000000010000",
42011 => "0000000000010000",42012 => "0000000000010000",
42013 => "0000000000010000",42014 => "0000000000010000",
42015 => "0000000000010000",42016 => "0000000000010000",
42017 => "0000000000010000",42018 => "0000000000010000",
42019 => "0000000000010000",42020 => "0000000000010000",
42021 => "0000000000010000",42022 => "0000000000010000",
42023 => "0000000000010000",42024 => "0000000000010000",
42025 => "0000000000010000",42026 => "0000000000010000",
42027 => "0000000000010000",42028 => "0000000000010000",
42029 => "0000000000010000",42030 => "0000000000010000",
42031 => "0000000000010000",42032 => "0000000000010000",
42033 => "0000000000010000",42034 => "0000000000010000",
42035 => "0000000000010000",42036 => "0000000000010000",
42037 => "0000000000010000",42038 => "0000000000010000",
42039 => "0000000000010000",42040 => "0000000000010000",
42041 => "0000000000010000",42042 => "0000000000010000",
42043 => "0000000000010000",42044 => "0000000000010000",
42045 => "0000000000010000",42046 => "0000000000010000",
42047 => "0000000000010000",42048 => "0000000000010000",
42049 => "0000000000010000",42050 => "0000000000010000",
42051 => "0000000000010000",42052 => "0000000000010000",
42053 => "0000000000010000",42054 => "0000000000010000",
42055 => "0000000000010000",42056 => "0000000000010000",
42057 => "0000000000010000",42058 => "0000000000010000",
42059 => "0000000000010000",42060 => "0000000000010000",
42061 => "0000000000010000",42062 => "0000000000010000",
42063 => "0000000000010000",42064 => "0000000000010000",
42065 => "0000000000010000",42066 => "0000000000010000",
42067 => "0000000000010000",42068 => "0000000000010000",
42069 => "0000000000010000",42070 => "0000000000010000",
42071 => "0000000000010000",42072 => "0000000000010000",
42073 => "0000000000010000",42074 => "0000000000010000",
42075 => "0000000000010000",42076 => "0000000000010000",
42077 => "0000000000010000",42078 => "0000000000010000",
42079 => "0000000000010000",42080 => "0000000000010000",
42081 => "0000000000010000",42082 => "0000000000010000",
42083 => "0000000000010000",42084 => "0000000000010000",
42085 => "0000000000010000",42086 => "0000000000010000",
42087 => "0000000000010000",42088 => "0000000000010000",
42089 => "0000000000010000",42090 => "0000000000010000",
42091 => "0000000000010000",42092 => "0000000000010000",
42093 => "0000000000010000",42094 => "0000000000010000",
42095 => "0000000000010000",42096 => "0000000000010000",
42097 => "0000000000010000",42098 => "0000000000010000",
42099 => "0000000000010000",42100 => "0000000000010000",
42101 => "0000000000010000",42102 => "0000000000010000",
42103 => "0000000000010000",42104 => "0000000000010000",
42105 => "0000000000010000",42106 => "0000000000010000",
42107 => "0000000000010000",42108 => "0000000000010000",
42109 => "0000000000010000",42110 => "0000000000010000",
42111 => "0000000000010000",42112 => "0000000000010000",
42113 => "0000000000010000",42114 => "0000000000010000",
42115 => "0000000000010000",42116 => "0000000000010000",
42117 => "0000000000010000",42118 => "0000000000010000",
42119 => "0000000000010000",42120 => "0000000000010000",
42121 => "0000000000010000",42122 => "0000000000010000",
42123 => "0000000000010000",42124 => "0000000000010000",
42125 => "0000000000010000",42126 => "0000000000010000",
42127 => "0000000000010000",42128 => "0000000000010000",
42129 => "0000000000010000",42130 => "0000000000010000",
42131 => "0000000000010000",42132 => "0000000000010000",
42133 => "0000000000010000",42134 => "0000000000010000",
42135 => "0000000000010000",42136 => "0000000000010000",
42137 => "0000000000010000",42138 => "0000000000010000",
42139 => "0000000000010000",42140 => "0000000000010000",
42141 => "0000000000010000",42142 => "0000000000010000",
42143 => "0000000000010000",42144 => "0000000000010000",
42145 => "0000000000010000",42146 => "0000000000010000",
42147 => "0000000000010000",42148 => "0000000000010000",
42149 => "0000000000010000",42150 => "0000000000010000",
42151 => "0000000000010000",42152 => "0000000000010000",
42153 => "0000000000010000",42154 => "0000000000010000",
42155 => "0000000000010000",42156 => "0000000000010000",
42157 => "0000000000010000",42158 => "0000000000010000",
42159 => "0000000000010000",42160 => "0000000000010000",
42161 => "0000000000010000",42162 => "0000000000010000",
42163 => "0000000000010000",42164 => "0000000000010000",
42165 => "0000000000010000",42166 => "0000000000010000",
42167 => "0000000000010000",42168 => "0000000000010000",
42169 => "0000000000010000",42170 => "0000000000010000",
42171 => "0000000000010000",42172 => "0000000000010000",
42173 => "0000000000010000",42174 => "0000000000010000",
42175 => "0000000000010000",42176 => "0000000000010000",
42177 => "0000000000010000",42178 => "0000000000010000",
42179 => "0000000000010000",42180 => "0000000000010000",
42181 => "0000000000010000",42182 => "0000000000010000",
42183 => "0000000000010000",42184 => "0000000000010000",
42185 => "0000000000010000",42186 => "0000000000010000",
42187 => "0000000000010000",42188 => "0000000000010000",
42189 => "0000000000010000",42190 => "0000000000010000",
42191 => "0000000000010000",42192 => "0000000000010000",
42193 => "0000000000010000",42194 => "0000000000010000",
42195 => "0000000000010000",42196 => "0000000000010000",
42197 => "0000000000010000",42198 => "0000000000010000",
42199 => "0000000000010000",42200 => "0000000000010000",
42201 => "0000000000010000",42202 => "0000000000010000",
42203 => "0000000000010000",42204 => "0000000000010000",
42205 => "0000000000010000",42206 => "0000000000010000",
42207 => "0000000000010000",42208 => "0000000000010000",
42209 => "0000000000010000",42210 => "0000000000010000",
42211 => "0000000000010000",42212 => "0000000000010000",
42213 => "0000000000010000",42214 => "0000000000010000",
42215 => "0000000000010000",42216 => "0000000000010000",
42217 => "0000000000010000",42218 => "0000000000010000",
42219 => "0000000000010000",42220 => "0000000000010000",
42221 => "0000000000010000",42222 => "0000000000010000",
42223 => "0000000000010000",42224 => "0000000000010000",
42225 => "0000000000010000",42226 => "0000000000010000",
42227 => "0000000000010000",42228 => "0000000000010000",
42229 => "0000000000010000",42230 => "0000000000010000",
42231 => "0000000000010000",42232 => "0000000000010000",
42233 => "0000000000010000",42234 => "0000000000010000",
42235 => "0000000000010000",42236 => "0000000000010000",
42237 => "0000000000010000",42238 => "0000000000010000",
42239 => "0000000000010000",42240 => "0000000000010000",
42241 => "0000000000010000",42242 => "0000000000010000",
42243 => "0000000000010000",42244 => "0000000000010000",
42245 => "0000000000010000",42246 => "0000000000010000",
42247 => "0000000000010000",42248 => "0000000000010000",
42249 => "0000000000010000",42250 => "0000000000010000",
42251 => "0000000000010000",42252 => "0000000000010000",
42253 => "0000000000010000",42254 => "0000000000010000",
42255 => "0000000000010000",42256 => "0000000000010000",
42257 => "0000000000010000",42258 => "0000000000010000",
42259 => "0000000000010000",42260 => "0000000000010000",
42261 => "0000000000010000",42262 => "0000000000010000",
42263 => "0000000000010000",42264 => "0000000000010000",
42265 => "0000000000010000",42266 => "0000000000010000",
42267 => "0000000000010000",42268 => "0000000000010000",
42269 => "0000000000010000",42270 => "0000000000010000",
42271 => "0000000000010000",42272 => "0000000000010000",
42273 => "0000000000010000",42274 => "0000000000010000",
42275 => "0000000000010000",42276 => "0000000000010000",
42277 => "0000000000010000",42278 => "0000000000010000",
42279 => "0000000000010000",42280 => "0000000000010000",
42281 => "0000000000010000",42282 => "0000000000010000",
42283 => "0000000000010000",42284 => "0000000000010000",
42285 => "0000000000010000",42286 => "0000000000010000",
42287 => "0000000000010000",42288 => "0000000000010000",
42289 => "0000000000010000",42290 => "0000000000010000",
42291 => "0000000000010000",42292 => "0000000000010000",
42293 => "0000000000010000",42294 => "0000000000010000",
42295 => "0000000000010000",42296 => "0000000000010000",
42297 => "0000000000010000",42298 => "0000000000010000",
42299 => "0000000000010000",42300 => "0000000000010000",
42301 => "0000000000010000",42302 => "0000000000010000",
42303 => "0000000000010000",42304 => "0000000000010000",
42305 => "0000000000010000",42306 => "0000000000010000",
42307 => "0000000000010000",42308 => "0000000000010000",
42309 => "0000000000010000",42310 => "0000000000010000",
42311 => "0000000000010000",42312 => "0000000000010000",
42313 => "0000000000010000",42314 => "0000000000010000",
42315 => "0000000000010000",42316 => "0000000000010000",
42317 => "0000000000010000",42318 => "0000000000010000",
42319 => "0000000000010000",42320 => "0000000000010000",
42321 => "0000000000010000",42322 => "0000000000010000",
42323 => "0000000000010000",42324 => "0000000000010000",
42325 => "0000000000010000",42326 => "0000000000010000",
42327 => "0000000000010000",42328 => "0000000000010000",
42329 => "0000000000010000",42330 => "0000000000010000",
42331 => "0000000000010000",42332 => "0000000000010000",
42333 => "0000000000010000",42334 => "0000000000010000",
42335 => "0000000000010000",42336 => "0000000000010000",
42337 => "0000000000010000",42338 => "0000000000010000",
42339 => "0000000000010000",42340 => "0000000000010000",
42341 => "0000000000010000",42342 => "0000000000010000",
42343 => "0000000000010000",42344 => "0000000000010000",
42345 => "0000000000010000",42346 => "0000000000010000",
42347 => "0000000000010000",42348 => "0000000000010000",
42349 => "0000000000010000",42350 => "0000000000010000",
42351 => "0000000000010000",42352 => "0000000000010000",
42353 => "0000000000010000",42354 => "0000000000010000",
42355 => "0000000000010000",42356 => "0000000000010000",
42357 => "0000000000010000",42358 => "0000000000010000",
42359 => "0000000000010000",42360 => "0000000000010000",
42361 => "0000000000010000",42362 => "0000000000010000",
42363 => "0000000000010000",42364 => "0000000000010000",
42365 => "0000000000010000",42366 => "0000000000010000",
42367 => "0000000000010000",42368 => "0000000000010000",
42369 => "0000000000010000",42370 => "0000000000010000",
42371 => "0000000000010000",42372 => "0000000000010000",
42373 => "0000000000010000",42374 => "0000000000010000",
42375 => "0000000000010000",42376 => "0000000000010000",
42377 => "0000000000010000",42378 => "0000000000010000",
42379 => "0000000000010000",42380 => "0000000000010000",
42381 => "0000000000010000",42382 => "0000000000010000",
42383 => "0000000000010000",42384 => "0000000000010000",
42385 => "0000000000010000",42386 => "0000000000010000",
42387 => "0000000000010000",42388 => "0000000000010000",
42389 => "0000000000010000",42390 => "0000000000010000",
42391 => "0000000000010000",42392 => "0000000000010000",
42393 => "0000000000010000",42394 => "0000000000010000",
42395 => "0000000000010000",42396 => "0000000000010000",
42397 => "0000000000010000",42398 => "0000000000010000",
42399 => "0000000000010000",42400 => "0000000000010000",
42401 => "0000000000010000",42402 => "0000000000010000",
42403 => "0000000000010000",42404 => "0000000000010000",
42405 => "0000000000010000",42406 => "0000000000010000",
42407 => "0000000000010000",42408 => "0000000000010000",
42409 => "0000000000010000",42410 => "0000000000010000",
42411 => "0000000000010000",42412 => "0000000000010000",
42413 => "0000000000010000",42414 => "0000000000010000",
42415 => "0000000000010000",42416 => "0000000000010000",
42417 => "0000000000010000",42418 => "0000000000010000",
42419 => "0000000000010000",42420 => "0000000000010000",
42421 => "0000000000010000",42422 => "0000000000010000",
42423 => "0000000000010000",42424 => "0000000000010000",
42425 => "0000000000010000",42426 => "0000000000010000",
42427 => "0000000000010000",42428 => "0000000000010000",
42429 => "0000000000010000",42430 => "0000000000010000",
42431 => "0000000000010000",42432 => "0000000000010000",
42433 => "0000000000010000",42434 => "0000000000010000",
42435 => "0000000000010000",42436 => "0000000000010000",
42437 => "0000000000010000",42438 => "0000000000010000",
42439 => "0000000000010000",42440 => "0000000000010000",
42441 => "0000000000010000",42442 => "0000000000010000",
42443 => "0000000000010000",42444 => "0000000000010000",
42445 => "0000000000010000",42446 => "0000000000010000",
42447 => "0000000000010000",42448 => "0000000000010000",
42449 => "0000000000010000",42450 => "0000000000010000",
42451 => "0000000000010000",42452 => "0000000000010000",
42453 => "0000000000010000",42454 => "0000000000010000",
42455 => "0000000000010000",42456 => "0000000000010000",
42457 => "0000000000010000",42458 => "0000000000010000",
42459 => "0000000000010000",42460 => "0000000000010000",
42461 => "0000000000010000",42462 => "0000000000010000",
42463 => "0000000000010000",42464 => "0000000000010000",
42465 => "0000000000010000",42466 => "0000000000010000",
42467 => "0000000000010000",42468 => "0000000000010000",
42469 => "0000000000010000",42470 => "0000000000010000",
42471 => "0000000000010000",42472 => "0000000000010000",
42473 => "0000000000010000",42474 => "0000000000010000",
42475 => "0000000000010000",42476 => "0000000000010000",
42477 => "0000000000010000",42478 => "0000000000010000",
42479 => "0000000000010000",42480 => "0000000000010000",
42481 => "0000000000010000",42482 => "0000000000010000",
42483 => "0000000000010000",42484 => "0000000000010000",
42485 => "0000000000010000",42486 => "0000000000010000",
42487 => "0000000000010000",42488 => "0000000000010000",
42489 => "0000000000010000",42490 => "0000000000010000",
42491 => "0000000000010000",42492 => "0000000000010000",
42493 => "0000000000010000",42494 => "0000000000010000",
42495 => "0000000000010000",42496 => "0000000000010000",
42497 => "0000000000010000",42498 => "0000000000010000",
42499 => "0000000000010000",42500 => "0000000000010000",
42501 => "0000000000010000",42502 => "0000000000010000",
42503 => "0000000000010000",42504 => "0000000000010000",
42505 => "0000000000010000",42506 => "0000000000010000",
42507 => "0000000000010000",42508 => "0000000000010000",
42509 => "0000000000010000",42510 => "0000000000010000",
42511 => "0000000000010000",42512 => "0000000000010000",
42513 => "0000000000010000",42514 => "0000000000010000",
42515 => "0000000000010000",42516 => "0000000000010000",
42517 => "0000000000010000",42518 => "0000000000010000",
42519 => "0000000000010000",42520 => "0000000000010000",
42521 => "0000000000010000",42522 => "0000000000010000",
42523 => "0000000000010000",42524 => "0000000000010000",
42525 => "0000000000010000",42526 => "0000000000010000",
42527 => "0000000000010000",42528 => "0000000000010000",
42529 => "0000000000010000",42530 => "0000000000010000",
42531 => "0000000000010000",42532 => "0000000000010000",
42533 => "0000000000010000",42534 => "0000000000010000",
42535 => "0000000000010000",42536 => "0000000000010000",
42537 => "0000000000010000",42538 => "0000000000010000",
42539 => "0000000000010000",42540 => "0000000000010000",
42541 => "0000000000010000",42542 => "0000000000010000",
42543 => "0000000000010000",42544 => "0000000000010000",
42545 => "0000000000010000",42546 => "0000000000010000",
42547 => "0000000000010000",42548 => "0000000000010000",
42549 => "0000000000010000",42550 => "0000000000010000",
42551 => "0000000000010000",42552 => "0000000000010000",
42553 => "0000000000010000",42554 => "0000000000010000",
42555 => "0000000000010000",42556 => "0000000000010000",
42557 => "0000000000010000",42558 => "0000000000010000",
42559 => "0000000000010000",42560 => "0000000000010000",
42561 => "0000000000010000",42562 => "0000000000010000",
42563 => "0000000000010000",42564 => "0000000000010000",
42565 => "0000000000010000",42566 => "0000000000010000",
42567 => "0000000000010000",42568 => "0000000000010000",
42569 => "0000000000010000",42570 => "0000000000010000",
42571 => "0000000000010000",42572 => "0000000000010000",
42573 => "0000000000010000",42574 => "0000000000010000",
42575 => "0000000000010000",42576 => "0000000000010000",
42577 => "0000000000010000",42578 => "0000000000010000",
42579 => "0000000000010000",42580 => "0000000000010000",
42581 => "0000000000010000",42582 => "0000000000010000",
42583 => "0000000000010000",42584 => "0000000000010000",
42585 => "0000000000010000",42586 => "0000000000010000",
42587 => "0000000000010000",42588 => "0000000000010000",
42589 => "0000000000010000",42590 => "0000000000010000",
42591 => "0000000000010000",42592 => "0000000000010000",
42593 => "0000000000010000",42594 => "0000000000010000",
42595 => "0000000000010000",42596 => "0000000000010000",
42597 => "0000000000010000",42598 => "0000000000010000",
42599 => "0000000000010000",42600 => "0000000000010000",
42601 => "0000000000010000",42602 => "0000000000010000",
42603 => "0000000000010000",42604 => "0000000000010000",
42605 => "0000000000010000",42606 => "0000000000010000",
42607 => "0000000000010000",42608 => "0000000000010000",
42609 => "0000000000010000",42610 => "0000000000010000",
42611 => "0000000000010000",42612 => "0000000000010000",
42613 => "0000000000010000",42614 => "0000000000010000",
42615 => "0000000000010000",42616 => "0000000000010000",
42617 => "0000000000010000",42618 => "0000000000010000",
42619 => "0000000000010000",42620 => "0000000000010000",
42621 => "0000000000010000",42622 => "0000000000010000",
42623 => "0000000000010000",42624 => "0000000000010000",
42625 => "0000000000010000",42626 => "0000000000010000",
42627 => "0000000000010000",42628 => "0000000000010000",
42629 => "0000000000010000",42630 => "0000000000001111",
42631 => "0000000000001111",42632 => "0000000000001111",
42633 => "0000000000001111",42634 => "0000000000001111",
42635 => "0000000000001111",42636 => "0000000000001111",
42637 => "0000000000001111",42638 => "0000000000001111",
42639 => "0000000000001111",42640 => "0000000000001111",
42641 => "0000000000001111",42642 => "0000000000001111",
42643 => "0000000000001111",42644 => "0000000000001111",
42645 => "0000000000001111",42646 => "0000000000001111",
42647 => "0000000000001111",42648 => "0000000000001111",
42649 => "0000000000001111",42650 => "0000000000001111",
42651 => "0000000000001111",42652 => "0000000000001111",
42653 => "0000000000001111",42654 => "0000000000001111",
42655 => "0000000000001111",42656 => "0000000000001111",
42657 => "0000000000001111",42658 => "0000000000001111",
42659 => "0000000000001111",42660 => "0000000000001111",
42661 => "0000000000001111",42662 => "0000000000001111",
42663 => "0000000000001111",42664 => "0000000000001111",
42665 => "0000000000001111",42666 => "0000000000001111",
42667 => "0000000000001111",42668 => "0000000000001111",
42669 => "0000000000001111",42670 => "0000000000001111",
42671 => "0000000000001111",42672 => "0000000000001111",
42673 => "0000000000001111",42674 => "0000000000001111",
42675 => "0000000000001111",42676 => "0000000000001111",
42677 => "0000000000001111",42678 => "0000000000001111",
42679 => "0000000000001111",42680 => "0000000000001111",
42681 => "0000000000001111",42682 => "0000000000001111",
42683 => "0000000000001111",42684 => "0000000000001111",
42685 => "0000000000001111",42686 => "0000000000001111",
42687 => "0000000000001111",42688 => "0000000000001111",
42689 => "0000000000001111",42690 => "0000000000001111",
42691 => "0000000000001111",42692 => "0000000000001111",
42693 => "0000000000001111",42694 => "0000000000001111",
42695 => "0000000000001111",42696 => "0000000000001111",
42697 => "0000000000001111",42698 => "0000000000001111",
42699 => "0000000000001111",42700 => "0000000000001111",
42701 => "0000000000001111",42702 => "0000000000001111",
42703 => "0000000000001111",42704 => "0000000000001111",
42705 => "0000000000001111",42706 => "0000000000001111",
42707 => "0000000000001111",42708 => "0000000000001111",
42709 => "0000000000001111",42710 => "0000000000001111",
42711 => "0000000000001111",42712 => "0000000000001111",
42713 => "0000000000001111",42714 => "0000000000001111",
42715 => "0000000000001111",42716 => "0000000000001111",
42717 => "0000000000001111",42718 => "0000000000001111",
42719 => "0000000000001111",42720 => "0000000000001111",
42721 => "0000000000001111",42722 => "0000000000001111",
42723 => "0000000000001111",42724 => "0000000000001111",
42725 => "0000000000001111",42726 => "0000000000001111",
42727 => "0000000000001111",42728 => "0000000000001111",
42729 => "0000000000001111",42730 => "0000000000001111",
42731 => "0000000000001111",42732 => "0000000000001111",
42733 => "0000000000001111",42734 => "0000000000001111",
42735 => "0000000000001111",42736 => "0000000000001111",
42737 => "0000000000001111",42738 => "0000000000001111",
42739 => "0000000000001111",42740 => "0000000000001111",
42741 => "0000000000001111",42742 => "0000000000001111",
42743 => "0000000000001111",42744 => "0000000000001111",
42745 => "0000000000001111",42746 => "0000000000001111",
42747 => "0000000000001111",42748 => "0000000000001111",
42749 => "0000000000001111",42750 => "0000000000001111",
42751 => "0000000000001111",42752 => "0000000000001111",
42753 => "0000000000001111",42754 => "0000000000001111",
42755 => "0000000000001111",42756 => "0000000000001111",
42757 => "0000000000001111",42758 => "0000000000001111",
42759 => "0000000000001111",42760 => "0000000000001111",
42761 => "0000000000001111",42762 => "0000000000001111",
42763 => "0000000000001111",42764 => "0000000000001111",
42765 => "0000000000001111",42766 => "0000000000001111",
42767 => "0000000000001111",42768 => "0000000000001111",
42769 => "0000000000001111",42770 => "0000000000001111",
42771 => "0000000000001111",42772 => "0000000000001111",
42773 => "0000000000001111",42774 => "0000000000001111",
42775 => "0000000000001111",42776 => "0000000000001111",
42777 => "0000000000001111",42778 => "0000000000001111",
42779 => "0000000000001111",42780 => "0000000000001111",
42781 => "0000000000001111",42782 => "0000000000001111",
42783 => "0000000000001111",42784 => "0000000000001111",
42785 => "0000000000001111",42786 => "0000000000001111",
42787 => "0000000000001111",42788 => "0000000000001111",
42789 => "0000000000001111",42790 => "0000000000001111",
42791 => "0000000000001111",42792 => "0000000000001111",
42793 => "0000000000001111",42794 => "0000000000001111",
42795 => "0000000000001111",42796 => "0000000000001111",
42797 => "0000000000001111",42798 => "0000000000001111",
42799 => "0000000000001111",42800 => "0000000000001111",
42801 => "0000000000001111",42802 => "0000000000001111",
42803 => "0000000000001111",42804 => "0000000000001111",
42805 => "0000000000001111",42806 => "0000000000001111",
42807 => "0000000000001111",42808 => "0000000000001111",
42809 => "0000000000001111",42810 => "0000000000001111",
42811 => "0000000000001111",42812 => "0000000000001111",
42813 => "0000000000001111",42814 => "0000000000001111",
42815 => "0000000000001111",42816 => "0000000000001111",
42817 => "0000000000001111",42818 => "0000000000001111",
42819 => "0000000000001111",42820 => "0000000000001111",
42821 => "0000000000001111",42822 => "0000000000001111",
42823 => "0000000000001111",42824 => "0000000000001111",
42825 => "0000000000001111",42826 => "0000000000001111",
42827 => "0000000000001111",42828 => "0000000000001111",
42829 => "0000000000001111",42830 => "0000000000001111",
42831 => "0000000000001111",42832 => "0000000000001111",
42833 => "0000000000001111",42834 => "0000000000001111",
42835 => "0000000000001111",42836 => "0000000000001111",
42837 => "0000000000001111",42838 => "0000000000001111",
42839 => "0000000000001111",42840 => "0000000000001111",
42841 => "0000000000001111",42842 => "0000000000001111",
42843 => "0000000000001111",42844 => "0000000000001111",
42845 => "0000000000001111",42846 => "0000000000001111",
42847 => "0000000000001111",42848 => "0000000000001111",
42849 => "0000000000001111",42850 => "0000000000001111",
42851 => "0000000000001111",42852 => "0000000000001111",
42853 => "0000000000001111",42854 => "0000000000001111",
42855 => "0000000000001111",42856 => "0000000000001111",
42857 => "0000000000001111",42858 => "0000000000001111",
42859 => "0000000000001111",42860 => "0000000000001111",
42861 => "0000000000001111",42862 => "0000000000001111",
42863 => "0000000000001111",42864 => "0000000000001111",
42865 => "0000000000001111",42866 => "0000000000001111",
42867 => "0000000000001111",42868 => "0000000000001111",
42869 => "0000000000001111",42870 => "0000000000001111",
42871 => "0000000000001111",42872 => "0000000000001111",
42873 => "0000000000001111",42874 => "0000000000001111",
42875 => "0000000000001111",42876 => "0000000000001111",
42877 => "0000000000001111",42878 => "0000000000001111",
42879 => "0000000000001111",42880 => "0000000000001111",
42881 => "0000000000001111",42882 => "0000000000001111",
42883 => "0000000000001111",42884 => "0000000000001111",
42885 => "0000000000001111",42886 => "0000000000001111",
42887 => "0000000000001111",42888 => "0000000000001111",
42889 => "0000000000001111",42890 => "0000000000001111",
42891 => "0000000000001111",42892 => "0000000000001111",
42893 => "0000000000001111",42894 => "0000000000001111",
42895 => "0000000000001111",42896 => "0000000000001111",
42897 => "0000000000001111",42898 => "0000000000001111",
42899 => "0000000000001111",42900 => "0000000000001111",
42901 => "0000000000001111",42902 => "0000000000001111",
42903 => "0000000000001111",42904 => "0000000000001111",
42905 => "0000000000001111",42906 => "0000000000001111",
42907 => "0000000000001111",42908 => "0000000000001111",
42909 => "0000000000001111",42910 => "0000000000001111",
42911 => "0000000000001111",42912 => "0000000000001111",
42913 => "0000000000001111",42914 => "0000000000001111",
42915 => "0000000000001111",42916 => "0000000000001111",
42917 => "0000000000001111",42918 => "0000000000001111",
42919 => "0000000000001111",42920 => "0000000000001111",
42921 => "0000000000001111",42922 => "0000000000001111",
42923 => "0000000000001111",42924 => "0000000000001111",
42925 => "0000000000001111",42926 => "0000000000001111",
42927 => "0000000000001111",42928 => "0000000000001111",
42929 => "0000000000001111",42930 => "0000000000001111",
42931 => "0000000000001111",42932 => "0000000000001111",
42933 => "0000000000001111",42934 => "0000000000001111",
42935 => "0000000000001111",42936 => "0000000000001111",
42937 => "0000000000001111",42938 => "0000000000001111",
42939 => "0000000000001111",42940 => "0000000000001111",
42941 => "0000000000001111",42942 => "0000000000001111",
42943 => "0000000000001111",42944 => "0000000000001111",
42945 => "0000000000001111",42946 => "0000000000001111",
42947 => "0000000000001111",42948 => "0000000000001111",
42949 => "0000000000001111",42950 => "0000000000001111",
42951 => "0000000000001111",42952 => "0000000000001111",
42953 => "0000000000001111",42954 => "0000000000001111",
42955 => "0000000000001111",42956 => "0000000000001111",
42957 => "0000000000001111",42958 => "0000000000001111",
42959 => "0000000000001111",42960 => "0000000000001111",
42961 => "0000000000001111",42962 => "0000000000001111",
42963 => "0000000000001111",42964 => "0000000000001111",
42965 => "0000000000001111",42966 => "0000000000001111",
42967 => "0000000000001111",42968 => "0000000000001111",
42969 => "0000000000001111",42970 => "0000000000001111",
42971 => "0000000000001111",42972 => "0000000000001111",
42973 => "0000000000001111",42974 => "0000000000001111",
42975 => "0000000000001111",42976 => "0000000000001111",
42977 => "0000000000001111",42978 => "0000000000001111",
42979 => "0000000000001111",42980 => "0000000000001111",
42981 => "0000000000001111",42982 => "0000000000001111",
42983 => "0000000000001111",42984 => "0000000000001111",
42985 => "0000000000001111",42986 => "0000000000001111",
42987 => "0000000000001111",42988 => "0000000000001111",
42989 => "0000000000001111",42990 => "0000000000001111",
42991 => "0000000000001111",42992 => "0000000000001111",
42993 => "0000000000001111",42994 => "0000000000001111",
42995 => "0000000000001111",42996 => "0000000000001111",
42997 => "0000000000001111",42998 => "0000000000001111",
42999 => "0000000000001111",43000 => "0000000000001111",
43001 => "0000000000001111",43002 => "0000000000001111",
43003 => "0000000000001111",43004 => "0000000000001111",
43005 => "0000000000001111",43006 => "0000000000001111",
43007 => "0000000000001111",43008 => "0000000000000111",
43009 => "0000000000000110",43010 => "0000000000000110",
43011 => "0000000000000101",43012 => "0000000000000101",
43013 => "0000000000000100",43014 => "0000000000000100",
43015 => "0000000000000011",43016 => "0000000000000011",
43017 => "0000000000000011",43018 => "0000000000000110",
43019 => "0000000000000110",43020 => "0000000000000110",
43021 => "0000000000000110",43022 => "0000000000000110",
43023 => "0000000000000110",43024 => "0000000000000110",
43025 => "0000000000000110",43026 => "0000000000000110",
43027 => "0000000000000110",43028 => "0000000000000110",
43029 => "0000000000000101",43030 => "0000000000000101",
43031 => "0000000000000101",43032 => "0000000000000101",
43033 => "0000000000000101",43034 => "0000000000000101",
43035 => "0000000000000101",43036 => "0000000000000101",
43037 => "0000000000000101",43038 => "0000000000000101",
43039 => "0000000000000101",43040 => "0000000000000101",
43041 => "0000000000000101",43042 => "0000000000000101",
43043 => "0000000000000101",43044 => "0000000000000101",
43045 => "0000000000000101",43046 => "0000000000000101",
43047 => "0000000000000101",43048 => "0000000000000101",
43049 => "0000000000000100",43050 => "0000000000000100",
43051 => "0000000000000100",43052 => "0000000000000100",
43053 => "0000000000000100",43054 => "0000000000000100",
43055 => "0000000000000100",43056 => "0000000000000100",
43057 => "0000000000000100",43058 => "0000000000000100",
43059 => "0000000000000100",43060 => "0000000000000100",
43061 => "0000000000000100",43062 => "0000000000000100",
43063 => "0000000000000100",43064 => "0000000000000100",
43065 => "0000000000000100",43066 => "0000000000000100",
43067 => "0000000000000100",43068 => "0000000000000100",
43069 => "0000000000000100",43070 => "0000000000000100",
43071 => "0000000000000100",43072 => "0000000000000100",
43073 => "0000000000000100",43074 => "0000000000000011",
43075 => "0000000000000011",43076 => "0000000000000011",
43077 => "0000000000000011",43078 => "0000000000000011",
43079 => "0000000000000011",43080 => "0000000000000011",
43081 => "0000000000000011",43082 => "0000000000000011",
43083 => "0000000000000011",43084 => "0000000000000011",
43085 => "0000000000000011",43086 => "0000000000000011",
43087 => "0000000000000011",43088 => "0000000000000011",
43089 => "0000000000000011",43090 => "0000000000000011",
43091 => "0000000000000011",43092 => "0000000000000011",
43093 => "0000000000000011",43094 => "0000000000000011",
43095 => "0000000000000011",43096 => "0000000000000011",
43097 => "0000000000000011",43098 => "0000000000000011",
43099 => "0000000000000011",43100 => "0000000000000011",
43101 => "0000000000000011",43102 => "0000000000000011",
43103 => "0000000000000011",43104 => "0000000000000011",
43105 => "0000000000000011",43106 => "0000000000000011",
43107 => "0000000000000011",43108 => "0000000000000110",
43109 => "0000000000000110",43110 => "0000000000000110",
43111 => "0000000000000110",43112 => "0000000000000110",
43113 => "0000000000000110",43114 => "0000000000000110",
43115 => "0000000000000110",43116 => "0000000000000110",
43117 => "0000000000000110",43118 => "0000000000000110",
43119 => "0000000000000110",43120 => "0000000000000110",
43121 => "0000000000000110",43122 => "0000000000000110",
43123 => "0000000000000110",43124 => "0000000000000110",
43125 => "0000000000000110",43126 => "0000000000000110",
43127 => "0000000000000110",43128 => "0000000000000110",
43129 => "0000000000000110",43130 => "0000000000000110",
43131 => "0000000000000110",43132 => "0000000000000110",
43133 => "0000000000000110",43134 => "0000000000000110",
43135 => "0000000000000110",43136 => "0000000000000110",
43137 => "0000000000000110",43138 => "0000000000000110",
43139 => "0000000000000110",43140 => "0000000000000110",
43141 => "0000000000000110",43142 => "0000000000000110",
43143 => "0000000000000110",43144 => "0000000000000110",
43145 => "0000000000000110",43146 => "0000000000000110",
43147 => "0000000000000110",43148 => "0000000000000110",
43149 => "0000000000000110",43150 => "0000000000000110",
43151 => "0000000000000110",43152 => "0000000000000110",
43153 => "0000000000000110",43154 => "0000000000000110",
43155 => "0000000000000110",43156 => "0000000000000110",
43157 => "0000000000000110",43158 => "0000000000000110",
43159 => "0000000000000110",43160 => "0000000000000110",
43161 => "0000000000000110",43162 => "0000000000000110",
43163 => "0000000000000110",43164 => "0000000000000110",
43165 => "0000000000000110",43166 => "0000000000000110",
43167 => "0000000000000110",43168 => "0000000000000110",
43169 => "0000000000000110",43170 => "0000000000000110",
43171 => "0000000000000110",43172 => "0000000000000110",
43173 => "0000000000000110",43174 => "0000000000000110",
43175 => "0000000000000110",43176 => "0000000000000110",
43177 => "0000000000000110",43178 => "0000000000000110",
43179 => "0000000000000110",43180 => "0000000000000110",
43181 => "0000000000000110",43182 => "0000000000000110",
43183 => "0000000000000110",43184 => "0000000000000110",
43185 => "0000000000000110",43186 => "0000000000000110",
43187 => "0000000000000110",43188 => "0000000000000110",
43189 => "0000000000000110",43190 => "0000000000000110",
43191 => "0000000000000110",43192 => "0000000000000110",
43193 => "0000000000000110",43194 => "0000000000000110",
43195 => "0000000000000110",43196 => "0000000000000110",
43197 => "0000000000000110",43198 => "0000000000000110",
43199 => "0000000000000110",43200 => "0000000000000110",
43201 => "0000000000000110",43202 => "0000000000000110",
43203 => "0000000000000110",43204 => "0000000000000110",
43205 => "0000000000000110",43206 => "0000000000000110",
43207 => "0000000000000110",43208 => "0000000000000110",
43209 => "0000000000000110",43210 => "0000000000000110",
43211 => "0000000000000110",43212 => "0000000000000101",
43213 => "0000000000000101",43214 => "0000000000000101",
43215 => "0000000000000101",43216 => "0000000000000101",
43217 => "0000000000000101",43218 => "0000000000000101",
43219 => "0000000000000101",43220 => "0000000000000101",
43221 => "0000000000000101",43222 => "0000000000000101",
43223 => "0000000000000101",43224 => "0000000000000101",
43225 => "0000000000000101",43226 => "0000000000000101",
43227 => "0000000000000101",43228 => "0000000000000101",
43229 => "0000000000000101",43230 => "0000000000000101",
43231 => "0000000000000101",43232 => "0000000000000101",
43233 => "0000000000000101",43234 => "0000000000000101",
43235 => "0000000000000101",43236 => "0000000000000101",
43237 => "0000000000000101",43238 => "0000000000000101",
43239 => "0000000000000101",43240 => "0000000000000101",
43241 => "0000000000000101",43242 => "0000000000000101",
43243 => "0000000000000101",43244 => "0000000000000101",
43245 => "0000000000000101",43246 => "0000000000000101",
43247 => "0000000000000101",43248 => "0000000000000101",
43249 => "0000000000000101",43250 => "0000000000000101",
43251 => "0000000000000101",43252 => "0000000000000101",
43253 => "0000000000000101",43254 => "0000000000000101",
43255 => "0000000000000101",43256 => "0000000000000101",
43257 => "0000000000000101",43258 => "0000000000000101",
43259 => "0000000000000101",43260 => "0000000000000101",
43261 => "0000000000000101",43262 => "0000000000000101",
43263 => "0000000000000101",43264 => "0000000000000101",
43265 => "0000000000000101",43266 => "0000000000000101",
43267 => "0000000000000101",43268 => "0000000000000101",
43269 => "0000000000000101",43270 => "0000000000000101",
43271 => "0000000000000101",43272 => "0000000000000101",
43273 => "0000000000000101",43274 => "0000000000000101",
43275 => "0000000000000101",43276 => "0000000000000101",
43277 => "0000000000000101",43278 => "0000000000000101",
43279 => "0000000000000101",43280 => "0000000000000101",
43281 => "0000000000000101",43282 => "0000000000000101",
43283 => "0000000000000101",43284 => "0000000000000101",
43285 => "0000000000000101",43286 => "0000000000000101",
43287 => "0000000000000101",43288 => "0000000000000101",
43289 => "0000000000000101",43290 => "0000000000000101",
43291 => "0000000000000101",43292 => "0000000000000101",
43293 => "0000000000000101",43294 => "0000000000000101",
43295 => "0000000000000101",43296 => "0000000000000101",
43297 => "0000000000000101",43298 => "0000000000000101",
43299 => "0000000000000101",43300 => "0000000000000101",
43301 => "0000000000000101",43302 => "0000000000000101",
43303 => "0000000000000101",43304 => "0000000000000101",
43305 => "0000000000000101",43306 => "0000000000000101",
43307 => "0000000000000101",43308 => "0000000000000101",
43309 => "0000000000000101",43310 => "0000000000000101",
43311 => "0000000000000101",43312 => "0000000000000101",
43313 => "0000000000000101",43314 => "0000000000000101",
43315 => "0000000000000101",43316 => "0000000000000101",
43317 => "0000000000000101",43318 => "0000000000000101",
43319 => "0000000000000101",43320 => "0000000000000101",
43321 => "0000000000000101",43322 => "0000000000000101",
43323 => "0000000000000101",43324 => "0000000000000101",
43325 => "0000000000000101",43326 => "0000000000000101",
43327 => "0000000000000101",43328 => "0000000000000101",
43329 => "0000000000000101",43330 => "0000000000000101",
43331 => "0000000000000101",43332 => "0000000000000101",
43333 => "0000000000000101",43334 => "0000000000000101",
43335 => "0000000000000101",43336 => "0000000000000101",
43337 => "0000000000000101",43338 => "0000000000000101",
43339 => "0000000000000101",43340 => "0000000000000101",
43341 => "0000000000000101",43342 => "0000000000000101",
43343 => "0000000000000101",43344 => "0000000000000101",
43345 => "0000000000000101",43346 => "0000000000000101",
43347 => "0000000000000101",43348 => "0000000000000101",
43349 => "0000000000000101",43350 => "0000000000000101",
43351 => "0000000000000101",43352 => "0000000000000101",
43353 => "0000000000000101",43354 => "0000000000000101",
43355 => "0000000000000101",43356 => "0000000000000101",
43357 => "0000000000000101",43358 => "0000000000000101",
43359 => "0000000000000101",43360 => "0000000000000101",
43361 => "0000000000000101",43362 => "0000000000000101",
43363 => "0000000000000101",43364 => "0000000000000101",
43365 => "0000000000000101",43366 => "0000000000000101",
43367 => "0000000000000101",43368 => "0000000000000101",
43369 => "0000000000000101",43370 => "0000000000000101",
43371 => "0000000000000101",43372 => "0000000000000101",
43373 => "0000000000000101",43374 => "0000000000000101",
43375 => "0000000000000101",43376 => "0000000000000101",
43377 => "0000000000000101",43378 => "0000000000000101",
43379 => "0000000000000101",43380 => "0000000000000101",
43381 => "0000000000000101",43382 => "0000000000000101",
43383 => "0000000000000101",43384 => "0000000000000101",
43385 => "0000000000000101",43386 => "0000000000000101",
43387 => "0000000000000101",43388 => "0000000000000101",
43389 => "0000000000000101",43390 => "0000000000000101",
43391 => "0000000000000101",43392 => "0000000000000101",
43393 => "0000000000000101",43394 => "0000000000000101",
43395 => "0000000000000101",43396 => "0000000000000101",
43397 => "0000000000000101",43398 => "0000000000000101",
43399 => "0000000000000101",43400 => "0000000000000101",
43401 => "0000000000000101",43402 => "0000000000000101",
43403 => "0000000000000101",43404 => "0000000000000101",
43405 => "0000000000000101",43406 => "0000000000000101",
43407 => "0000000000000101",43408 => "0000000000000101",
43409 => "0000000000000101",43410 => "0000000000000101",
43411 => "0000000000000101",43412 => "0000000000000100",
43413 => "0000000000000100",43414 => "0000000000000100",
43415 => "0000000000000100",43416 => "0000000000000100",
43417 => "0000000000000100",43418 => "0000000000000100",
43419 => "0000000000000100",43420 => "0000000000000100",
43421 => "0000000000000100",43422 => "0000000000000100",
43423 => "0000000000000100",43424 => "0000000000000100",
43425 => "0000000000000100",43426 => "0000000000000100",
43427 => "0000000000000100",43428 => "0000000000000100",
43429 => "0000000000000100",43430 => "0000000000000100",
43431 => "0000000000000100",43432 => "0000000000000100",
43433 => "0000000000000100",43434 => "0000000000000100",
43435 => "0000000000000100",43436 => "0000000000000100",
43437 => "0000000000000100",43438 => "0000000000000100",
43439 => "0000000000000100",43440 => "0000000000000100",
43441 => "0000000000000100",43442 => "0000000000000100",
43443 => "0000000000000100",43444 => "0000000000000100",
43445 => "0000000000000100",43446 => "0000000000000100",
43447 => "0000000000000100",43448 => "0000000000000100",
43449 => "0000000000000100",43450 => "0000000000000100",
43451 => "0000000000000100",43452 => "0000000000000100",
43453 => "0000000000000100",43454 => "0000000000000100",
43455 => "0000000000000100",43456 => "0000000000000100",
43457 => "0000000000000100",43458 => "0000000000000100",
43459 => "0000000000000100",43460 => "0000000000000100",
43461 => "0000000000000100",43462 => "0000000000000100",
43463 => "0000000000000100",43464 => "0000000000000100",
43465 => "0000000000000100",43466 => "0000000000000100",
43467 => "0000000000000100",43468 => "0000000000000100",
43469 => "0000000000000100",43470 => "0000000000000100",
43471 => "0000000000000100",43472 => "0000000000000100",
43473 => "0000000000000100",43474 => "0000000000000100",
43475 => "0000000000000100",43476 => "0000000000000100",
43477 => "0000000000000100",43478 => "0000000000000100",
43479 => "0000000000000100",43480 => "0000000000000100",
43481 => "0000000000000100",43482 => "0000000000000100",
43483 => "0000000000000100",43484 => "0000000000000100",
43485 => "0000000000000100",43486 => "0000000000000100",
43487 => "0000000000000100",43488 => "0000000000000100",
43489 => "0000000000000100",43490 => "0000000000000100",
43491 => "0000000000000100",43492 => "0000000000000100",
43493 => "0000000000000100",43494 => "0000000000000100",
43495 => "0000000000000100",43496 => "0000000000000100",
43497 => "0000000000000100",43498 => "0000000000000100",
43499 => "0000000000000100",43500 => "0000000000000100",
43501 => "0000000000000100",43502 => "0000000000000100",
43503 => "0000000000000100",43504 => "0000000000000100",
43505 => "0000000000000100",43506 => "0000000000000100",
43507 => "0000000000000100",43508 => "0000000000000100",
43509 => "0000000000000100",43510 => "0000000000000100",
43511 => "0000000000000100",43512 => "0000000000000100",
43513 => "0000000000000100",43514 => "0000000000000100",
43515 => "0000000000000100",43516 => "0000000000000100",
43517 => "0000000000000100",43518 => "0000000000000100",
43519 => "0000000000000100",43520 => "0000000000000100",
43521 => "0000000000000100",43522 => "0000000000000100",
43523 => "0000000000000100",43524 => "0000000000000100",
43525 => "0000000000000100",43526 => "0000000000000100",
43527 => "0000000000000100",43528 => "0000000000000100",
43529 => "0000000000000100",43530 => "0000000000000100",
43531 => "0000000000000100",43532 => "0000000000000100",
43533 => "0000000000000100",43534 => "0000000000000100",
43535 => "0000000000000100",43536 => "0000000000000100",
43537 => "0000000000000100",43538 => "0000000000000100",
43539 => "0000000000000100",43540 => "0000000000000100",
43541 => "0000000000000100",43542 => "0000000000000100",
43543 => "0000000000000100",43544 => "0000000000000100",
43545 => "0000000000000100",43546 => "0000000000000100",
43547 => "0000000000000100",43548 => "0000000000000100",
43549 => "0000000000000100",43550 => "0000000000000100",
43551 => "0000000000000100",43552 => "0000000000000100",
43553 => "0000000000000100",43554 => "0000000000000100",
43555 => "0000000000000100",43556 => "0000000000000100",
43557 => "0000000000000100",43558 => "0000000000000100",
43559 => "0000000000000100",43560 => "0000000000000100",
43561 => "0000000000000100",43562 => "0000000000000100",
43563 => "0000000000000100",43564 => "0000000000000100",
43565 => "0000000000000100",43566 => "0000000000000100",
43567 => "0000000000000100",43568 => "0000000000000100",
43569 => "0000000000000100",43570 => "0000000000000100",
43571 => "0000000000000100",43572 => "0000000000000100",
43573 => "0000000000000100",43574 => "0000000000000100",
43575 => "0000000000000100",43576 => "0000000000000100",
43577 => "0000000000000100",43578 => "0000000000000100",
43579 => "0000000000000100",43580 => "0000000000000100",
43581 => "0000000000000100",43582 => "0000000000000100",
43583 => "0000000000000100",43584 => "0000000000000100",
43585 => "0000000000000100",43586 => "0000000000000100",
43587 => "0000000000000100",43588 => "0000000000000100",
43589 => "0000000000000100",43590 => "0000000000000100",
43591 => "0000000000000100",43592 => "0000000000000100",
43593 => "0000000000000100",43594 => "0000000000000100",
43595 => "0000000000000100",43596 => "0000000000000100",
43597 => "0000000000000100",43598 => "0000000000000100",
43599 => "0000000000000100",43600 => "0000000000000100",
43601 => "0000000000000100",43602 => "0000000000000100",
43603 => "0000000000000100",43604 => "0000000000000100",
43605 => "0000000000000100",43606 => "0000000000000100",
43607 => "0000000000000100",43608 => "0000000000000100",
43609 => "0000000000000100",43610 => "0000000000000100",
43611 => "0000000000000100",43612 => "0000000000000100",
43613 => "0000000000000100",43614 => "0000000000000100",
43615 => "0000000000000100",43616 => "0000000000000100",
43617 => "0000000000000100",43618 => "0000000000000100",
43619 => "0000000000000100",43620 => "0000000000000100",
43621 => "0000000000000100",43622 => "0000000000000100",
43623 => "0000000000000100",43624 => "0000000000000100",
43625 => "0000000000000100",43626 => "0000000000000100",
43627 => "0000000000000100",43628 => "0000000000000100",
43629 => "0000000000000100",43630 => "0000000000000100",
43631 => "0000000000000100",43632 => "0000000000000100",
43633 => "0000000000000100",43634 => "0000000000000100",
43635 => "0000000000000100",43636 => "0000000000000100",
43637 => "0000000000000100",43638 => "0000000000000100",
43639 => "0000000000000100",43640 => "0000000000000100",
43641 => "0000000000000100",43642 => "0000000000000100",
43643 => "0000000000000100",43644 => "0000000000000100",
43645 => "0000000000000100",43646 => "0000000000000100",
43647 => "0000000000000100",43648 => "0000000000000100",
43649 => "0000000000000100",43650 => "0000000000000100",
43651 => "0000000000000100",43652 => "0000000000000100",
43653 => "0000000000000100",43654 => "0000000000000100",
43655 => "0000000000000100",43656 => "0000000000000100",
43657 => "0000000000000100",43658 => "0000000000000100",
43659 => "0000000000000100",43660 => "0000000000000100",
43661 => "0000000000000100",43662 => "0000000000000100",
43663 => "0000000000000011",43664 => "0000000000000011",
43665 => "0000000000000011",43666 => "0000000000000011",
43667 => "0000000000000011",43668 => "0000000000000011",
43669 => "0000000000000011",43670 => "0000000000000011",
43671 => "0000000000000011",43672 => "0000000000000011",
43673 => "0000000000000011",43674 => "0000000000000011",
43675 => "0000000000000011",43676 => "0000000000000011",
43677 => "0000000000000011",43678 => "0000000000000011",
43679 => "0000000000000011",43680 => "0000000000000011",
43681 => "0000000000000011",43682 => "0000000000000011",
43683 => "0000000000000011",43684 => "0000000000000011",
43685 => "0000000000000011",43686 => "0000000000000011",
43687 => "0000000000000011",43688 => "0000000000000011",
43689 => "0000000000000011",43690 => "0000000000000011",
43691 => "0000000000000011",43692 => "0000000000000011",
43693 => "0000000000000011",43694 => "0000000000000011",
43695 => "0000000000000011",43696 => "0000000000000011",
43697 => "0000000000000011",43698 => "0000000000000011",
43699 => "0000000000000011",43700 => "0000000000000011",
43701 => "0000000000000011",43702 => "0000000000000011",
43703 => "0000000000000011",43704 => "0000000000000011",
43705 => "0000000000000011",43706 => "0000000000000011",
43707 => "0000000000000011",43708 => "0000000000000011",
43709 => "0000000000000011",43710 => "0000000000000011",
43711 => "0000000000000011",43712 => "0000000000000011",
43713 => "0000000000000011",43714 => "0000000000000011",
43715 => "0000000000000011",43716 => "0000000000000011",
43717 => "0000000000000011",43718 => "0000000000000011",
43719 => "0000000000000011",43720 => "0000000000000011",
43721 => "0000000000000011",43722 => "0000000000000011",
43723 => "0000000000000011",43724 => "0000000000000011",
43725 => "0000000000000011",43726 => "0000000000000011",
43727 => "0000000000000011",43728 => "0000000000000011",
43729 => "0000000000000011",43730 => "0000000000000011",
43731 => "0000000000000011",43732 => "0000000000000011",
43733 => "0000000000000011",43734 => "0000000000000011",
43735 => "0000000000000011",43736 => "0000000000000011",
43737 => "0000000000000011",43738 => "0000000000000011",
43739 => "0000000000000011",43740 => "0000000000000011",
43741 => "0000000000000011",43742 => "0000000000000011",
43743 => "0000000000000011",43744 => "0000000000000011",
43745 => "0000000000000011",43746 => "0000000000000011",
43747 => "0000000000000011",43748 => "0000000000000011",
43749 => "0000000000000011",43750 => "0000000000000011",
43751 => "0000000000000011",43752 => "0000000000000011",
43753 => "0000000000000011",43754 => "0000000000000011",
43755 => "0000000000000011",43756 => "0000000000000011",
43757 => "0000000000000011",43758 => "0000000000000011",
43759 => "0000000000000011",43760 => "0000000000000011",
43761 => "0000000000000011",43762 => "0000000000000011",
43763 => "0000000000000011",43764 => "0000000000000011",
43765 => "0000000000000011",43766 => "0000000000000011",
43767 => "0000000000000011",43768 => "0000000000000011",
43769 => "0000000000000011",43770 => "0000000000000011",
43771 => "0000000000000011",43772 => "0000000000000011",
43773 => "0000000000000011",43774 => "0000000000000011",
43775 => "0000000000000011",43776 => "0000000000000011",
43777 => "0000000000000011",43778 => "0000000000000011",
43779 => "0000000000000011",43780 => "0000000000000011",
43781 => "0000000000000011",43782 => "0000000000000011",
43783 => "0000000000000011",43784 => "0000000000000011",
43785 => "0000000000000011",43786 => "0000000000000011",
43787 => "0000000000000011",43788 => "0000000000000011",
43789 => "0000000000000011",43790 => "0000000000000011",
43791 => "0000000000000011",43792 => "0000000000000011",
43793 => "0000000000000011",43794 => "0000000000000011",
43795 => "0000000000000011",43796 => "0000000000000011",
43797 => "0000000000000011",43798 => "0000000000000011",
43799 => "0000000000000011",43800 => "0000000000000011",
43801 => "0000000000000011",43802 => "0000000000000011",
43803 => "0000000000000011",43804 => "0000000000000011",
43805 => "0000000000000011",43806 => "0000000000000011",
43807 => "0000000000000011",43808 => "0000000000000011",
43809 => "0000000000000011",43810 => "0000000000000011",
43811 => "0000000000000011",43812 => "0000000000000011",
43813 => "0000000000000011",43814 => "0000000000000011",
43815 => "0000000000000011",43816 => "0000000000000011",
43817 => "0000000000000011",43818 => "0000000000000011",
43819 => "0000000000000011",43820 => "0000000000000011",
43821 => "0000000000000011",43822 => "0000000000000011",
43823 => "0000000000000011",43824 => "0000000000000011",
43825 => "0000000000000011",43826 => "0000000000000011",
43827 => "0000000000000011",43828 => "0000000000000011",
43829 => "0000000000000011",43830 => "0000000000000011",
43831 => "0000000000000011",43832 => "0000000000000011",
43833 => "0000000000000011",43834 => "0000000000000011",
43835 => "0000000000000011",43836 => "0000000000000011",
43837 => "0000000000000011",43838 => "0000000000000011",
43839 => "0000000000000011",43840 => "0000000000000011",
43841 => "0000000000000011",43842 => "0000000000000011",
43843 => "0000000000000011",43844 => "0000000000000011",
43845 => "0000000000000011",43846 => "0000000000000011",
43847 => "0000000000000011",43848 => "0000000000000011",
43849 => "0000000000000011",43850 => "0000000000000011",
43851 => "0000000000000011",43852 => "0000000000000011",
43853 => "0000000000000011",43854 => "0000000000000011",
43855 => "0000000000000011",43856 => "0000000000000011",
43857 => "0000000000000011",43858 => "0000000000000011",
43859 => "0000000000000011",43860 => "0000000000000011",
43861 => "0000000000000011",43862 => "0000000000000011",
43863 => "0000000000000011",43864 => "0000000000000011",
43865 => "0000000000000011",43866 => "0000000000000011",
43867 => "0000000000000011",43868 => "0000000000000011",
43869 => "0000000000000011",43870 => "0000000000000011",
43871 => "0000000000000011",43872 => "0000000000000011",
43873 => "0000000000000011",43874 => "0000000000000011",
43875 => "0000000000000011",43876 => "0000000000000011",
43877 => "0000000000000011",43878 => "0000000000000011",
43879 => "0000000000000011",43880 => "0000000000000011",
43881 => "0000000000000011",43882 => "0000000000000011",
43883 => "0000000000000011",43884 => "0000000000000011",
43885 => "0000000000000011",43886 => "0000000000000011",
43887 => "0000000000000011",43888 => "0000000000000011",
43889 => "0000000000000011",43890 => "0000000000000011",
43891 => "0000000000000011",43892 => "0000000000000011",
43893 => "0000000000000011",43894 => "0000000000000011",
43895 => "0000000000000011",43896 => "0000000000000011",
43897 => "0000000000000011",43898 => "0000000000000011",
43899 => "0000000000000011",43900 => "0000000000000011",
43901 => "0000000000000011",43902 => "0000000000000011",
43903 => "0000000000000011",43904 => "0000000000000011",
43905 => "0000000000000011",43906 => "0000000000000011",
43907 => "0000000000000011",43908 => "0000000000000011",
43909 => "0000000000000011",43910 => "0000000000000011",
43911 => "0000000000000011",43912 => "0000000000000011",
43913 => "0000000000000011",43914 => "0000000000000011",
43915 => "0000000000000011",43916 => "0000000000000011",
43917 => "0000000000000011",43918 => "0000000000000011",
43919 => "0000000000000011",43920 => "0000000000000011",
43921 => "0000000000000011",43922 => "0000000000000011",
43923 => "0000000000000011",43924 => "0000000000000011",
43925 => "0000000000000011",43926 => "0000000000000011",
43927 => "0000000000000011",43928 => "0000000000000011",
43929 => "0000000000000011",43930 => "0000000000000011",
43931 => "0000000000000011",43932 => "0000000000000011",
43933 => "0000000000000011",43934 => "0000000000000011",
43935 => "0000000000000011",43936 => "0000000000000011",
43937 => "0000000000000011",43938 => "0000000000000011",
43939 => "0000000000000011",43940 => "0000000000000011",
43941 => "0000000000000011",43942 => "0000000000000011",
43943 => "0000000000000011",43944 => "0000000000000011",
43945 => "0000000000000011",43946 => "0000000000000011",
43947 => "0000000000000011",43948 => "0000000000000011",
43949 => "0000000000000011",43950 => "0000000000000011",
43951 => "0000000000000011",43952 => "0000000000000011",
43953 => "0000000000000011",43954 => "0000000000000011",
43955 => "0000000000000011",43956 => "0000000000000011",
43957 => "0000000000000011",43958 => "0000000000000011",
43959 => "0000000000000011",43960 => "0000000000000011",
43961 => "0000000000000011",43962 => "0000000000000011",
43963 => "0000000000000011",43964 => "0000000000000011",
43965 => "0000000000000011",43966 => "0000000000000011",
43967 => "0000000000000011",43968 => "0000000000000011",
43969 => "0000000000000011",43970 => "0000000000000011",
43971 => "0000000000000011",43972 => "0000000000000011",
43973 => "0000000000000011",43974 => "0000000000000011",
43975 => "0000000000000011",43976 => "0000000000000011",
43977 => "0000000000000011",43978 => "0000000000000011",
43979 => "0000000000000011",43980 => "0000000000000011",
43981 => "0000000000000011",43982 => "0000000000000011",
43983 => "0000000000000011",43984 => "0000000000000011",
43985 => "0000000000000011",43986 => "0000000000000011",
43987 => "0000000000000011",43988 => "0000000000000011",
43989 => "0000000000000011",43990 => "0000000000000011",
43991 => "0000000000000011",43992 => "0000000000000011",
43993 => "0000000000000011",43994 => "0000000000000011",
43995 => "0000000000000011",43996 => "0000000000000011",
43997 => "0000000000000011",43998 => "0000000000000011",
43999 => "0000000000000011",44000 => "0000000000000010",
44001 => "0000000000000010",44002 => "0000000000000010",
44003 => "0000000000000010",44004 => "0000000000000010",
44005 => "0000000000000010",44006 => "0000000000000010",
44007 => "0000000000000010",44008 => "0000000000000110",
44009 => "0000000000000110",44010 => "0000000000000110",
44011 => "0000000000000110",44012 => "0000000000000110",
44013 => "0000000000000110",44014 => "0000000000000110",
44015 => "0000000000000110",44016 => "0000000000000110",
44017 => "0000000000000110",44018 => "0000000000000110",
44019 => "0000000000000110",44020 => "0000000000000110",
44021 => "0000000000000110",44022 => "0000000000000110",
44023 => "0000000000000110",44024 => "0000000000000110",
44025 => "0000000000000110",44026 => "0000000000000110",
44027 => "0000000000000110",44028 => "0000000000000110",
44029 => "0000000000000110",44030 => "0000000000000110",
44031 => "0000000000000110",44032 => "0000000000000110",
44033 => "0000000000000110",44034 => "0000000000000110",
44035 => "0000000000000110",44036 => "0000000000000110",
44037 => "0000000000000110",44038 => "0000000000000110",
44039 => "0000000000000110",44040 => "0000000000000110",
44041 => "0000000000000110",44042 => "0000000000000110",
44043 => "0000000000000110",44044 => "0000000000000110",
44045 => "0000000000000110",44046 => "0000000000000110",
44047 => "0000000000000110",44048 => "0000000000000110",
44049 => "0000000000000110",44050 => "0000000000000110",
44051 => "0000000000000110",44052 => "0000000000000110",
44053 => "0000000000000110",44054 => "0000000000000110",
44055 => "0000000000000110",44056 => "0000000000000110",
44057 => "0000000000000110",44058 => "0000000000000110",
44059 => "0000000000000110",44060 => "0000000000000110",
44061 => "0000000000000110",44062 => "0000000000000110",
44063 => "0000000000000110",44064 => "0000000000000110",
44065 => "0000000000000110",44066 => "0000000000000110",
44067 => "0000000000000110",44068 => "0000000000000110",
44069 => "0000000000000110",44070 => "0000000000000110",
44071 => "0000000000000110",44072 => "0000000000000110",
44073 => "0000000000000110",44074 => "0000000000000110",
44075 => "0000000000000110",44076 => "0000000000000110",
44077 => "0000000000000110",44078 => "0000000000000110",
44079 => "0000000000000110",44080 => "0000000000000110",
44081 => "0000000000000110",44082 => "0000000000000110",
44083 => "0000000000000110",44084 => "0000000000000110",
44085 => "0000000000000110",44086 => "0000000000000110",
44087 => "0000000000000110",44088 => "0000000000000110",
44089 => "0000000000000110",44090 => "0000000000000110",
44091 => "0000000000000110",44092 => "0000000000000110",
44093 => "0000000000000110",44094 => "0000000000000110",
44095 => "0000000000000110",44096 => "0000000000000110",
44097 => "0000000000000110",44098 => "0000000000000110",
44099 => "0000000000000110",44100 => "0000000000000110",
44101 => "0000000000000110",44102 => "0000000000000110",
44103 => "0000000000000110",44104 => "0000000000000110",
44105 => "0000000000000110",44106 => "0000000000000110",
44107 => "0000000000000110",44108 => "0000000000000110",
44109 => "0000000000000110",44110 => "0000000000000110",
44111 => "0000000000000110",44112 => "0000000000000110",
44113 => "0000000000000110",44114 => "0000000000000110",
44115 => "0000000000000110",44116 => "0000000000000110",
44117 => "0000000000000110",44118 => "0000000000000110",
44119 => "0000000000000110",44120 => "0000000000000110",
44121 => "0000000000000110",44122 => "0000000000000110",
44123 => "0000000000000110",44124 => "0000000000000110",
44125 => "0000000000000110",44126 => "0000000000000110",
44127 => "0000000000000110",44128 => "0000000000000110",
44129 => "0000000000000110",44130 => "0000000000000110",
44131 => "0000000000000110",44132 => "0000000000000110",
44133 => "0000000000000110",44134 => "0000000000000110",
44135 => "0000000000000110",44136 => "0000000000000110",
44137 => "0000000000000110",44138 => "0000000000000110",
44139 => "0000000000000110",44140 => "0000000000000110",
44141 => "0000000000000110",44142 => "0000000000000110",
44143 => "0000000000000110",44144 => "0000000000000110",
44145 => "0000000000000110",44146 => "0000000000000110",
44147 => "0000000000000110",44148 => "0000000000000110",
44149 => "0000000000000110",44150 => "0000000000000110",
44151 => "0000000000000110",44152 => "0000000000000110",
44153 => "0000000000000110",44154 => "0000000000000110",
44155 => "0000000000000110",44156 => "0000000000000110",
44157 => "0000000000000110",44158 => "0000000000000110",
44159 => "0000000000000110",44160 => "0000000000000110",
44161 => "0000000000000110",44162 => "0000000000000110",
44163 => "0000000000000110",44164 => "0000000000000110",
44165 => "0000000000000110",44166 => "0000000000000110",
44167 => "0000000000000110",44168 => "0000000000000110",
44169 => "0000000000000110",44170 => "0000000000000110",
44171 => "0000000000000110",44172 => "0000000000000110",
44173 => "0000000000000110",44174 => "0000000000000110",
44175 => "0000000000000110",44176 => "0000000000000110",
44177 => "0000000000000110",44178 => "0000000000000110",
44179 => "0000000000000110",44180 => "0000000000000110",
44181 => "0000000000000110",44182 => "0000000000000110",
44183 => "0000000000000110",44184 => "0000000000000110",
44185 => "0000000000000110",44186 => "0000000000000110",
44187 => "0000000000000110",44188 => "0000000000000110",
44189 => "0000000000000110",44190 => "0000000000000110",
44191 => "0000000000000110",44192 => "0000000000000110",
44193 => "0000000000000110",44194 => "0000000000000110",
44195 => "0000000000000110",44196 => "0000000000000110",
44197 => "0000000000000110",44198 => "0000000000000110",
44199 => "0000000000000110",44200 => "0000000000000110",
44201 => "0000000000000110",44202 => "0000000000000110",
44203 => "0000000000000110",44204 => "0000000000000110",
44205 => "0000000000000110",44206 => "0000000000000110",
44207 => "0000000000000110",44208 => "0000000000000110",
44209 => "0000000000000110",44210 => "0000000000000110",
44211 => "0000000000000110",44212 => "0000000000000110",
44213 => "0000000000000110",44214 => "0000000000000110",
44215 => "0000000000000110",44216 => "0000000000000110",
44217 => "0000000000000110",44218 => "0000000000000110",
44219 => "0000000000000110",44220 => "0000000000000110",
44221 => "0000000000000110",44222 => "0000000000000110",
44223 => "0000000000000110",44224 => "0000000000000110",
44225 => "0000000000000110",44226 => "0000000000000110",
44227 => "0000000000000110",44228 => "0000000000000110",
44229 => "0000000000000110",44230 => "0000000000000110",
44231 => "0000000000000110",44232 => "0000000000000110",
44233 => "0000000000000110",44234 => "0000000000000110",
44235 => "0000000000000110",44236 => "0000000000000110",
44237 => "0000000000000110",44238 => "0000000000000110",
44239 => "0000000000000110",44240 => "0000000000000110",
44241 => "0000000000000110",44242 => "0000000000000110",
44243 => "0000000000000110",44244 => "0000000000000110",
44245 => "0000000000000110",44246 => "0000000000000110",
44247 => "0000000000000110",44248 => "0000000000000110",
44249 => "0000000000000110",44250 => "0000000000000110",
44251 => "0000000000000110",44252 => "0000000000000110",
44253 => "0000000000000110",44254 => "0000000000000110",
44255 => "0000000000000110",44256 => "0000000000000110",
44257 => "0000000000000110",44258 => "0000000000000110",
44259 => "0000000000000110",44260 => "0000000000000110",
44261 => "0000000000000110",44262 => "0000000000000110",
44263 => "0000000000000110",44264 => "0000000000000110",
44265 => "0000000000000110",44266 => "0000000000000110",
44267 => "0000000000000110",44268 => "0000000000000110",
44269 => "0000000000000110",44270 => "0000000000000110",
44271 => "0000000000000110",44272 => "0000000000000110",
44273 => "0000000000000110",44274 => "0000000000000110",
44275 => "0000000000000110",44276 => "0000000000000110",
44277 => "0000000000000110",44278 => "0000000000000110",
44279 => "0000000000000110",44280 => "0000000000000110",
44281 => "0000000000000110",44282 => "0000000000000110",
44283 => "0000000000000110",44284 => "0000000000000110",
44285 => "0000000000000110",44286 => "0000000000000110",
44287 => "0000000000000110",44288 => "0000000000000110",
44289 => "0000000000000110",44290 => "0000000000000110",
44291 => "0000000000000110",44292 => "0000000000000110",
44293 => "0000000000000110",44294 => "0000000000000110",
44295 => "0000000000000110",44296 => "0000000000000110",
44297 => "0000000000000110",44298 => "0000000000000110",
44299 => "0000000000000110",44300 => "0000000000000110",
44301 => "0000000000000110",44302 => "0000000000000110",
44303 => "0000000000000110",44304 => "0000000000000110",
44305 => "0000000000000110",44306 => "0000000000000110",
44307 => "0000000000000110",44308 => "0000000000000110",
44309 => "0000000000000110",44310 => "0000000000000110",
44311 => "0000000000000110",44312 => "0000000000000110",
44313 => "0000000000000110",44314 => "0000000000000110",
44315 => "0000000000000110",44316 => "0000000000000110",
44317 => "0000000000000110",44318 => "0000000000000110",
44319 => "0000000000000110",44320 => "0000000000000110",
44321 => "0000000000000110",44322 => "0000000000000110",
44323 => "0000000000000110",44324 => "0000000000000110",
44325 => "0000000000000110",44326 => "0000000000000110",
44327 => "0000000000000110",44328 => "0000000000000110",
44329 => "0000000000000110",44330 => "0000000000000110",
44331 => "0000000000000110",44332 => "0000000000000110",
44333 => "0000000000000110",44334 => "0000000000000110",
44335 => "0000000000000110",44336 => "0000000000000110",
44337 => "0000000000000110",44338 => "0000000000000110",
44339 => "0000000000000110",44340 => "0000000000000110",
44341 => "0000000000000110",44342 => "0000000000000110",
44343 => "0000000000000110",44344 => "0000000000000110",
44345 => "0000000000000110",44346 => "0000000000000110",
44347 => "0000000000000110",44348 => "0000000000000110",
44349 => "0000000000000110",44350 => "0000000000000110",
44351 => "0000000000000110",44352 => "0000000000000110",
44353 => "0000000000000110",44354 => "0000000000000110",
44355 => "0000000000000110",44356 => "0000000000000110",
44357 => "0000000000000110",44358 => "0000000000000110",
44359 => "0000000000000110",44360 => "0000000000000110",
44361 => "0000000000000110",44362 => "0000000000000110",
44363 => "0000000000000110",44364 => "0000000000000110",
44365 => "0000000000000110",44366 => "0000000000000110",
44367 => "0000000000000110",44368 => "0000000000000110",
44369 => "0000000000000110",44370 => "0000000000000110",
44371 => "0000000000000110",44372 => "0000000000000110",
44373 => "0000000000000110",44374 => "0000000000000110",
44375 => "0000000000000110",44376 => "0000000000000110",
44377 => "0000000000000110",44378 => "0000000000000110",
44379 => "0000000000000110",44380 => "0000000000000110",
44381 => "0000000000000110",44382 => "0000000000000110",
44383 => "0000000000000110",44384 => "0000000000000110",
44385 => "0000000000000110",44386 => "0000000000000110",
44387 => "0000000000000110",44388 => "0000000000000110",
44389 => "0000000000000110",44390 => "0000000000000110",
44391 => "0000000000000110",44392 => "0000000000000110",
44393 => "0000000000000110",44394 => "0000000000000110",
44395 => "0000000000000110",44396 => "0000000000000110",
44397 => "0000000000000110",44398 => "0000000000000110",
44399 => "0000000000000110",44400 => "0000000000000110",
44401 => "0000000000000110",44402 => "0000000000000110",
44403 => "0000000000000110",44404 => "0000000000000110",
44405 => "0000000000000110",44406 => "0000000000000110",
44407 => "0000000000000110",44408 => "0000000000000110",
44409 => "0000000000000110",44410 => "0000000000000110",
44411 => "0000000000000110",44412 => "0000000000000110",
44413 => "0000000000000110",44414 => "0000000000000110",
44415 => "0000000000000110",44416 => "0000000000000110",
44417 => "0000000000000110",44418 => "0000000000000110",
44419 => "0000000000000110",44420 => "0000000000000110",
44421 => "0000000000000110",44422 => "0000000000000110",
44423 => "0000000000000110",44424 => "0000000000000110",
44425 => "0000000000000110",44426 => "0000000000000110",
44427 => "0000000000000110",44428 => "0000000000000110",
44429 => "0000000000000110",44430 => "0000000000000110",
44431 => "0000000000000110",44432 => "0000000000000110",
44433 => "0000000000000110",44434 => "0000000000000110",
44435 => "0000000000000110",44436 => "0000000000000110",
44437 => "0000000000000110",44438 => "0000000000000110",
44439 => "0000000000000110",44440 => "0000000000000110",
44441 => "0000000000000110",44442 => "0000000000000110",
44443 => "0000000000000110",44444 => "0000000000000110",
44445 => "0000000000000110",44446 => "0000000000000110",
44447 => "0000000000000110",44448 => "0000000000000110",
44449 => "0000000000000110",44450 => "0000000000000110",
44451 => "0000000000000110",44452 => "0000000000000110",
44453 => "0000000000000110",44454 => "0000000000000110",
44455 => "0000000000000110",44456 => "0000000000000110",
44457 => "0000000000000110",44458 => "0000000000000110",
44459 => "0000000000000110",44460 => "0000000000000110",
44461 => "0000000000000110",44462 => "0000000000000110",
44463 => "0000000000000110",44464 => "0000000000000110",
44465 => "0000000000000110",44466 => "0000000000000110",
44467 => "0000000000000110",44468 => "0000000000000110",
44469 => "0000000000000110",44470 => "0000000000000110",
44471 => "0000000000000110",44472 => "0000000000000110",
44473 => "0000000000000110",44474 => "0000000000000110",
44475 => "0000000000000110",44476 => "0000000000000110",
44477 => "0000000000000110",44478 => "0000000000000110",
44479 => "0000000000000110",44480 => "0000000000000110",
44481 => "0000000000000110",44482 => "0000000000000110",
44483 => "0000000000000110",44484 => "0000000000000110",
44485 => "0000000000000110",44486 => "0000000000000110",
44487 => "0000000000000110",44488 => "0000000000000110",
44489 => "0000000000000110",44490 => "0000000000000110",
44491 => "0000000000000110",44492 => "0000000000000110",
44493 => "0000000000000110",44494 => "0000000000000110",
44495 => "0000000000000110",44496 => "0000000000000110",
44497 => "0000000000000110",44498 => "0000000000000110",
44499 => "0000000000000110",44500 => "0000000000000110",
44501 => "0000000000000110",44502 => "0000000000000110",
44503 => "0000000000000110",44504 => "0000000000000110",
44505 => "0000000000000110",44506 => "0000000000000110",
44507 => "0000000000000110",44508 => "0000000000000110",
44509 => "0000000000000110",44510 => "0000000000000110",
44511 => "0000000000000110",44512 => "0000000000000110",
44513 => "0000000000000110",44514 => "0000000000000110",
44515 => "0000000000000110",44516 => "0000000000000110",
44517 => "0000000000000110",44518 => "0000000000000110",
44519 => "0000000000000110",44520 => "0000000000000110",
44521 => "0000000000000110",44522 => "0000000000000110",
44523 => "0000000000000110",44524 => "0000000000000110",
44525 => "0000000000000110",44526 => "0000000000000110",
44527 => "0000000000000110",44528 => "0000000000000110",
44529 => "0000000000000110",44530 => "0000000000000110",
44531 => "0000000000000110",44532 => "0000000000000110",
44533 => "0000000000000110",44534 => "0000000000000110",
44535 => "0000000000000110",44536 => "0000000000000110",
44537 => "0000000000000110",44538 => "0000000000000110",
44539 => "0000000000000110",44540 => "0000000000000110",
44541 => "0000000000000110",44542 => "0000000000000110",
44543 => "0000000000000110",44544 => "0000000000000110",
44545 => "0000000000000110",44546 => "0000000000000110",
44547 => "0000000000000110",44548 => "0000000000000110",
44549 => "0000000000000110",44550 => "0000000000000110",
44551 => "0000000000000110",44552 => "0000000000000110",
44553 => "0000000000000110",44554 => "0000000000000110",
44555 => "0000000000000110",44556 => "0000000000000110",
44557 => "0000000000000110",44558 => "0000000000000110",
44559 => "0000000000000110",44560 => "0000000000000110",
44561 => "0000000000000110",44562 => "0000000000000110",
44563 => "0000000000000110",44564 => "0000000000000110",
44565 => "0000000000000110",44566 => "0000000000000110",
44567 => "0000000000000110",44568 => "0000000000000110",
44569 => "0000000000000110",44570 => "0000000000000110",
44571 => "0000000000000110",44572 => "0000000000000110",
44573 => "0000000000000110",44574 => "0000000000000110",
44575 => "0000000000000110",44576 => "0000000000000110",
44577 => "0000000000000110",44578 => "0000000000000110",
44579 => "0000000000000110",44580 => "0000000000000110",
44581 => "0000000000000110",44582 => "0000000000000110",
44583 => "0000000000000110",44584 => "0000000000000110",
44585 => "0000000000000110",44586 => "0000000000000110",
44587 => "0000000000000110",44588 => "0000000000000110",
44589 => "0000000000000110",44590 => "0000000000000110",
44591 => "0000000000000110",44592 => "0000000000000110",
44593 => "0000000000000110",44594 => "0000000000000110",
44595 => "0000000000000110",44596 => "0000000000000110",
44597 => "0000000000000110",44598 => "0000000000000110",
44599 => "0000000000000110",44600 => "0000000000000110",
44601 => "0000000000000110",44602 => "0000000000000110",
44603 => "0000000000000110",44604 => "0000000000000110",
44605 => "0000000000000110",44606 => "0000000000000110",
44607 => "0000000000000110",44608 => "0000000000000110",
44609 => "0000000000000110",44610 => "0000000000000110",
44611 => "0000000000000110",44612 => "0000000000000110",
44613 => "0000000000000110",44614 => "0000000000000110",
44615 => "0000000000000110",44616 => "0000000000000110",
44617 => "0000000000000110",44618 => "0000000000000110",
44619 => "0000000000000110",44620 => "0000000000000110",
44621 => "0000000000000110",44622 => "0000000000000110",
44623 => "0000000000000110",44624 => "0000000000000110",
44625 => "0000000000000110",44626 => "0000000000000110",
44627 => "0000000000000110",44628 => "0000000000000110",
44629 => "0000000000000110",44630 => "0000000000000110",
44631 => "0000000000000110",44632 => "0000000000000110",
44633 => "0000000000000110",44634 => "0000000000000110",
44635 => "0000000000000110",44636 => "0000000000000110",
44637 => "0000000000000110",44638 => "0000000000000110",
44639 => "0000000000000110",44640 => "0000000000000110",
44641 => "0000000000000110",44642 => "0000000000000110",
44643 => "0000000000000110",44644 => "0000000000000110",
44645 => "0000000000000110",44646 => "0000000000000110",
44647 => "0000000000000110",44648 => "0000000000000110",
44649 => "0000000000000110",44650 => "0000000000000110",
44651 => "0000000000000110",44652 => "0000000000000110",
44653 => "0000000000000110",44654 => "0000000000000110",
44655 => "0000000000000110",44656 => "0000000000000110",
44657 => "0000000000000110",44658 => "0000000000000110",
44659 => "0000000000000110",44660 => "0000000000000110",
44661 => "0000000000000110",44662 => "0000000000000110",
44663 => "0000000000000110",44664 => "0000000000000110",
44665 => "0000000000000110",44666 => "0000000000000110",
44667 => "0000000000000110",44668 => "0000000000000110",
44669 => "0000000000000110",44670 => "0000000000000110",
44671 => "0000000000000110",44672 => "0000000000000110",
44673 => "0000000000000110",44674 => "0000000000000110",
44675 => "0000000000000110",44676 => "0000000000000110",
44677 => "0000000000000110",44678 => "0000000000000110",
44679 => "0000000000000110",44680 => "0000000000000110",
44681 => "0000000000000110",44682 => "0000000000000110",
44683 => "0000000000000110",44684 => "0000000000000110",
44685 => "0000000000000110",44686 => "0000000000000110",
44687 => "0000000000000110",44688 => "0000000000000110",
44689 => "0000000000000110",44690 => "0000000000000110",
44691 => "0000000000000110",44692 => "0000000000000110",
44693 => "0000000000000110",44694 => "0000000000000110",
44695 => "0000000000000110",44696 => "0000000000000110",
44697 => "0000000000000110",44698 => "0000000000000110",
44699 => "0000000000000110",44700 => "0000000000000110",
44701 => "0000000000000110",44702 => "0000000000000110",
44703 => "0000000000000110",44704 => "0000000000000110",
44705 => "0000000000000110",44706 => "0000000000000110",
44707 => "0000000000000110",44708 => "0000000000000110",
44709 => "0000000000000110",44710 => "0000000000000110",
44711 => "0000000000000110",44712 => "0000000000000110",
44713 => "0000000000000110",44714 => "0000000000000110",
44715 => "0000000000000110",44716 => "0000000000000110",
44717 => "0000000000000110",44718 => "0000000000000110",
44719 => "0000000000000110",44720 => "0000000000000110",
44721 => "0000000000000110",44722 => "0000000000000110",
44723 => "0000000000000110",44724 => "0000000000000110",
44725 => "0000000000000110",44726 => "0000000000000110",
44727 => "0000000000000110",44728 => "0000000000000110",
44729 => "0000000000000110",44730 => "0000000000000110",
44731 => "0000000000000110",44732 => "0000000000000110",
44733 => "0000000000000110",44734 => "0000000000000110",
44735 => "0000000000000110",44736 => "0000000000000110",
44737 => "0000000000000110",44738 => "0000000000000110",
44739 => "0000000000000110",44740 => "0000000000000110",
44741 => "0000000000000110",44742 => "0000000000000110",
44743 => "0000000000000110",44744 => "0000000000000110",
44745 => "0000000000000110",44746 => "0000000000000110",
44747 => "0000000000000110",44748 => "0000000000000110",
44749 => "0000000000000110",44750 => "0000000000000110",
44751 => "0000000000000110",44752 => "0000000000000110",
44753 => "0000000000000110",44754 => "0000000000000110",
44755 => "0000000000000110",44756 => "0000000000000110",
44757 => "0000000000000110",44758 => "0000000000000110",
44759 => "0000000000000110",44760 => "0000000000000110",
44761 => "0000000000000110",44762 => "0000000000000110",
44763 => "0000000000000110",44764 => "0000000000000110",
44765 => "0000000000000110",44766 => "0000000000000110",
44767 => "0000000000000110",44768 => "0000000000000110",
44769 => "0000000000000110",44770 => "0000000000000110",
44771 => "0000000000000110",44772 => "0000000000000110",
44773 => "0000000000000110",44774 => "0000000000000110",
44775 => "0000000000000110",44776 => "0000000000000110",
44777 => "0000000000000110",44778 => "0000000000000110",
44779 => "0000000000000110",44780 => "0000000000000110",
44781 => "0000000000000110",44782 => "0000000000000110",
44783 => "0000000000000110",44784 => "0000000000000110",
44785 => "0000000000000110",44786 => "0000000000000110",
44787 => "0000000000000110",44788 => "0000000000000110",
44789 => "0000000000000110",44790 => "0000000000000110",
44791 => "0000000000000110",44792 => "0000000000000110",
44793 => "0000000000000110",44794 => "0000000000000110",
44795 => "0000000000000110",44796 => "0000000000000110",
44797 => "0000000000000110",44798 => "0000000000000110",
44799 => "0000000000000110",44800 => "0000000000000110",
44801 => "0000000000000110",44802 => "0000000000000110",
44803 => "0000000000000110",44804 => "0000000000000110",
44805 => "0000000000000110",44806 => "0000000000000110",
44807 => "0000000000000110",44808 => "0000000000000110",
44809 => "0000000000000110",44810 => "0000000000000110",
44811 => "0000000000000110",44812 => "0000000000000110",
44813 => "0000000000000110",44814 => "0000000000000110",
44815 => "0000000000000110",44816 => "0000000000000110",
44817 => "0000000000000110",44818 => "0000000000000110",
44819 => "0000000000000110",44820 => "0000000000000110",
44821 => "0000000000000110",44822 => "0000000000000110",
44823 => "0000000000000110",44824 => "0000000000000110",
44825 => "0000000000000110",44826 => "0000000000000110",
44827 => "0000000000000110",44828 => "0000000000000110",
44829 => "0000000000000110",44830 => "0000000000000110",
44831 => "0000000000000110",44832 => "0000000000000110",
44833 => "0000000000000110",44834 => "0000000000000110",
44835 => "0000000000000110",44836 => "0000000000000110",
44837 => "0000000000000110",44838 => "0000000000000110",
44839 => "0000000000000110",44840 => "0000000000000110",
44841 => "0000000000000110",44842 => "0000000000000110",
44843 => "0000000000000110",44844 => "0000000000000110",
44845 => "0000000000000110",44846 => "0000000000000110",
44847 => "0000000000000110",44848 => "0000000000000110",
44849 => "0000000000000110",44850 => "0000000000000110",
44851 => "0000000000000110",44852 => "0000000000000110",
44853 => "0000000000000110",44854 => "0000000000000110",
44855 => "0000000000000110",44856 => "0000000000000110",
44857 => "0000000000000110",44858 => "0000000000000110",
44859 => "0000000000000110",44860 => "0000000000000110",
44861 => "0000000000000110",44862 => "0000000000000110",
44863 => "0000000000000110",44864 => "0000000000000110",
44865 => "0000000000000110",44866 => "0000000000000110",
44867 => "0000000000000110",44868 => "0000000000000110",
44869 => "0000000000000110",44870 => "0000000000000110",
44871 => "0000000000000110",44872 => "0000000000000110",
44873 => "0000000000000110",44874 => "0000000000000110",
44875 => "0000000000000110",44876 => "0000000000000110",
44877 => "0000000000000110",44878 => "0000000000000110",
44879 => "0000000000000110",44880 => "0000000000000110",
44881 => "0000000000000110",44882 => "0000000000000110",
44883 => "0000000000000110",44884 => "0000000000000110",
44885 => "0000000000000110",44886 => "0000000000000110",
44887 => "0000000000000110",44888 => "0000000000000110",
44889 => "0000000000000110",44890 => "0000000000000110",
44891 => "0000000000000110",44892 => "0000000000000110",
44893 => "0000000000000110",44894 => "0000000000000110",
44895 => "0000000000000110",44896 => "0000000000000110",
44897 => "0000000000000110",44898 => "0000000000000110",
44899 => "0000000000000110",44900 => "0000000000000110",
44901 => "0000000000000110",44902 => "0000000000000110",
44903 => "0000000000000110",44904 => "0000000000000110",
44905 => "0000000000000110",44906 => "0000000000000110",
44907 => "0000000000000110",44908 => "0000000000000110",
44909 => "0000000000000110",44910 => "0000000000000110",
44911 => "0000000000000110",44912 => "0000000000000110",
44913 => "0000000000000110",44914 => "0000000000000110",
44915 => "0000000000000110",44916 => "0000000000000110",
44917 => "0000000000000110",44918 => "0000000000000110",
44919 => "0000000000000110",44920 => "0000000000000110",
44921 => "0000000000000110",44922 => "0000000000000110",
44923 => "0000000000000110",44924 => "0000000000000110",
44925 => "0000000000000110",44926 => "0000000000000110",
44927 => "0000000000000110",44928 => "0000000000000110",
44929 => "0000000000000110",44930 => "0000000000000110",
44931 => "0000000000000110",44932 => "0000000000000110",
44933 => "0000000000000110",44934 => "0000000000000110",
44935 => "0000000000000110",44936 => "0000000000000110",
44937 => "0000000000000110",44938 => "0000000000000110",
44939 => "0000000000000110",44940 => "0000000000000110",
44941 => "0000000000000110",44942 => "0000000000000110",
44943 => "0000000000000110",44944 => "0000000000000110",
44945 => "0000000000000110",44946 => "0000000000000110",
44947 => "0000000000000110",44948 => "0000000000000110",
44949 => "0000000000000110",44950 => "0000000000000110",
44951 => "0000000000000110",44952 => "0000000000000110",
44953 => "0000000000000110",44954 => "0000000000000110",
44955 => "0000000000000110",44956 => "0000000000000110",
44957 => "0000000000000110",44958 => "0000000000000110",
44959 => "0000000000000110",44960 => "0000000000000110",
44961 => "0000000000000110",44962 => "0000000000000110",
44963 => "0000000000000110",44964 => "0000000000000110",
44965 => "0000000000000110",44966 => "0000000000000110",
44967 => "0000000000000110",44968 => "0000000000000110",
44969 => "0000000000000110",44970 => "0000000000000110",
44971 => "0000000000000110",44972 => "0000000000000110",
44973 => "0000000000000110",44974 => "0000000000000110",
44975 => "0000000000000110",44976 => "0000000000000110",
44977 => "0000000000000110",44978 => "0000000000000110",
44979 => "0000000000000110",44980 => "0000000000000110",
44981 => "0000000000000110",44982 => "0000000000000110",
44983 => "0000000000000110",44984 => "0000000000000110",
44985 => "0000000000000110",44986 => "0000000000000110",
44987 => "0000000000000110",44988 => "0000000000000110",
44989 => "0000000000000110",44990 => "0000000000000110",
44991 => "0000000000000110",44992 => "0000000000000110",
44993 => "0000000000000110",44994 => "0000000000000110",
44995 => "0000000000000110",44996 => "0000000000000110",
44997 => "0000000000000110",44998 => "0000000000000110",
44999 => "0000000000000110",45000 => "0000000000000110",
45001 => "0000000000000110",45002 => "0000000000000110",
45003 => "0000000000000110",45004 => "0000000000000110",
45005 => "0000000000000110",45006 => "0000000000000110",
45007 => "0000000000000110",45008 => "0000000000000110",
45009 => "0000000000000110",45010 => "0000000000000110",
45011 => "0000000000000110",45012 => "0000000000000110",
45013 => "0000000000000110",45014 => "0000000000000110",
45015 => "0000000000000110",45016 => "0000000000000110",
45017 => "0000000000000110",45018 => "0000000000000110",
45019 => "0000000000000110",45020 => "0000000000000110",
45021 => "0000000000000110",45022 => "0000000000000110",
45023 => "0000000000000110",45024 => "0000000000000110",
45025 => "0000000000000110",45026 => "0000000000000110",
45027 => "0000000000000110",45028 => "0000000000000110",
45029 => "0000000000000110",45030 => "0000000000000110",
45031 => "0000000000000110",45032 => "0000000000000110",
45033 => "0000000000000110",45034 => "0000000000000110",
45035 => "0000000000000110",45036 => "0000000000000110",
45037 => "0000000000000110",45038 => "0000000000000110",
45039 => "0000000000000101",45040 => "0000000000000101",
45041 => "0000000000000101",45042 => "0000000000000101",
45043 => "0000000000000101",45044 => "0000000000000101",
45045 => "0000000000000101",45046 => "0000000000000101",
45047 => "0000000000000101",45048 => "0000000000000101",
45049 => "0000000000000101",45050 => "0000000000000101",
45051 => "0000000000000101",45052 => "0000000000000101",
45053 => "0000000000000101",45054 => "0000000000000101",
45055 => "0000000000000101",45056 => "0000000000000010",
45057 => "0000000000000010",45058 => "0000000000000010",
45059 => "0000000000000010",45060 => "0000000000000010",
45061 => "0000000000000010",45062 => "0000000000000001",
45063 => "0000000000000001",45064 => "0000000000000001",
45065 => "0000000000000001",45066 => "0000000000000010",
45067 => "0000000000000010",45068 => "0000000000000010",
45069 => "0000000000000010",45070 => "0000000000000010",
45071 => "0000000000000010",45072 => "0000000000000010",
45073 => "0000000000000010",45074 => "0000000000000010",
45075 => "0000000000000010",45076 => "0000000000000010",
45077 => "0000000000000010",45078 => "0000000000000010",
45079 => "0000000000000010",45080 => "0000000000000010",
45081 => "0000000000000010",45082 => "0000000000000010",
45083 => "0000000000000010",45084 => "0000000000000010",
45085 => "0000000000000010",45086 => "0000000000000010",
45087 => "0000000000000010",45088 => "0000000000000010",
45089 => "0000000000000010",45090 => "0000000000000010",
45091 => "0000000000000010",45092 => "0000000000000010",
45093 => "0000000000000010",45094 => "0000000000000010",
45095 => "0000000000000010",45096 => "0000000000000010",
45097 => "0000000000000010",45098 => "0000000000000010",
45099 => "0000000000000010",45100 => "0000000000000010",
45101 => "0000000000000010",45102 => "0000000000000010",
45103 => "0000000000000010",45104 => "0000000000000010",
45105 => "0000000000000010",45106 => "0000000000000010",
45107 => "0000000000000001",45108 => "0000000000000001",
45109 => "0000000000000001",45110 => "0000000000000001",
45111 => "0000000000000001",45112 => "0000000000000001",
45113 => "0000000000000001",45114 => "0000000000000001",
45115 => "0000000000000001",45116 => "0000000000000001",
45117 => "0000000000000001",45118 => "0000000000000001",
45119 => "0000000000000001",45120 => "0000000000000001",
45121 => "0000000000000001",45122 => "0000000000000001",
45123 => "0000000000000001",45124 => "0000000000000001",
45125 => "0000000000000001",45126 => "0000000000000001",
45127 => "0000000000000001",45128 => "0000000000000001",
45129 => "0000000000000001",45130 => "0000000000000001",
45131 => "0000000000000001",45132 => "0000000000000001",
45133 => "0000000000000001",45134 => "0000000000000001",
45135 => "0000000000000001",45136 => "0000000000000001",
45137 => "0000000000000001",45138 => "0000000000000001",
45139 => "0000000000000001",45140 => "0000000000000001",
45141 => "0000000000000001",45142 => "0000000000000001",
45143 => "0000000000000001",45144 => "0000000000000001",
45145 => "0000000000000001",45146 => "0000000000000001",
45147 => "0000000000000001",45148 => "0000000000000001",
45149 => "0000000000000001",45150 => "0000000000000001",
45151 => "0000000000000001",45152 => "0000000000000001",
45153 => "0000000000000001",45154 => "0000000000000001",
45155 => "0000000000000001",45156 => "0000000000000010",
45157 => "0000000000000010",45158 => "0000000000000010",
45159 => "0000000000000010",45160 => "0000000000000010",
45161 => "0000000000000010",45162 => "0000000000000010",
45163 => "0000000000000010",45164 => "0000000000000010",
45165 => "0000000000000010",45166 => "0000000000000010",
45167 => "0000000000000010",45168 => "0000000000000010",
45169 => "0000000000000010",45170 => "0000000000000010",
45171 => "0000000000000010",45172 => "0000000000000010",
45173 => "0000000000000010",45174 => "0000000000000010",
45175 => "0000000000000010",45176 => "0000000000000010",
45177 => "0000000000000010",45178 => "0000000000000010",
45179 => "0000000000000010",45180 => "0000000000000010",
45181 => "0000000000000010",45182 => "0000000000000010",
45183 => "0000000000000010",45184 => "0000000000000010",
45185 => "0000000000000010",45186 => "0000000000000010",
45187 => "0000000000000010",45188 => "0000000000000010",
45189 => "0000000000000010",45190 => "0000000000000010",
45191 => "0000000000000010",45192 => "0000000000000010",
45193 => "0000000000000010",45194 => "0000000000000010",
45195 => "0000000000000010",45196 => "0000000000000010",
45197 => "0000000000000010",45198 => "0000000000000010",
45199 => "0000000000000010",45200 => "0000000000000010",
45201 => "0000000000000010",45202 => "0000000000000010",
45203 => "0000000000000010",45204 => "0000000000000010",
45205 => "0000000000000010",45206 => "0000000000000010",
45207 => "0000000000000010",45208 => "0000000000000010",
45209 => "0000000000000010",45210 => "0000000000000010",
45211 => "0000000000000010",45212 => "0000000000000010",
45213 => "0000000000000010",45214 => "0000000000000010",
45215 => "0000000000000010",45216 => "0000000000000010",
45217 => "0000000000000010",45218 => "0000000000000010",
45219 => "0000000000000010",45220 => "0000000000000010",
45221 => "0000000000000010",45222 => "0000000000000010",
45223 => "0000000000000010",45224 => "0000000000000010",
45225 => "0000000000000010",45226 => "0000000000000010",
45227 => "0000000000000010",45228 => "0000000000000010",
45229 => "0000000000000010",45230 => "0000000000000010",
45231 => "0000000000000010",45232 => "0000000000000010",
45233 => "0000000000000010",45234 => "0000000000000010",
45235 => "0000000000000010",45236 => "0000000000000010",
45237 => "0000000000000010",45238 => "0000000000000010",
45239 => "0000000000000010",45240 => "0000000000000010",
45241 => "0000000000000010",45242 => "0000000000000010",
45243 => "0000000000000010",45244 => "0000000000000010",
45245 => "0000000000000010",45246 => "0000000000000010",
45247 => "0000000000000010",45248 => "0000000000000010",
45249 => "0000000000000010",45250 => "0000000000000010",
45251 => "0000000000000010",45252 => "0000000000000010",
45253 => "0000000000000010",45254 => "0000000000000010",
45255 => "0000000000000010",45256 => "0000000000000010",
45257 => "0000000000000010",45258 => "0000000000000010",
45259 => "0000000000000010",45260 => "0000000000000010",
45261 => "0000000000000010",45262 => "0000000000000010",
45263 => "0000000000000010",45264 => "0000000000000010",
45265 => "0000000000000010",45266 => "0000000000000010",
45267 => "0000000000000010",45268 => "0000000000000010",
45269 => "0000000000000010",45270 => "0000000000000010",
45271 => "0000000000000010",45272 => "0000000000000010",
45273 => "0000000000000010",45274 => "0000000000000010",
45275 => "0000000000000010",45276 => "0000000000000010",
45277 => "0000000000000010",45278 => "0000000000000010",
45279 => "0000000000000010",45280 => "0000000000000010",
45281 => "0000000000000010",45282 => "0000000000000010",
45283 => "0000000000000010",45284 => "0000000000000010",
45285 => "0000000000000010",45286 => "0000000000000010",
45287 => "0000000000000010",45288 => "0000000000000010",
45289 => "0000000000000010",45290 => "0000000000000010",
45291 => "0000000000000010",45292 => "0000000000000010",
45293 => "0000000000000010",45294 => "0000000000000010",
45295 => "0000000000000010",45296 => "0000000000000010",
45297 => "0000000000000010",45298 => "0000000000000010",
45299 => "0000000000000010",45300 => "0000000000000010",
45301 => "0000000000000010",45302 => "0000000000000010",
45303 => "0000000000000010",45304 => "0000000000000010",
45305 => "0000000000000010",45306 => "0000000000000010",
45307 => "0000000000000010",45308 => "0000000000000010",
45309 => "0000000000000010",45310 => "0000000000000010",
45311 => "0000000000000010",45312 => "0000000000000010",
45313 => "0000000000000010",45314 => "0000000000000010",
45315 => "0000000000000010",45316 => "0000000000000010",
45317 => "0000000000000010",45318 => "0000000000000010",
45319 => "0000000000000010",45320 => "0000000000000010",
45321 => "0000000000000010",45322 => "0000000000000010",
45323 => "0000000000000010",45324 => "0000000000000010",
45325 => "0000000000000010",45326 => "0000000000000010",
45327 => "0000000000000010",45328 => "0000000000000010",
45329 => "0000000000000010",45330 => "0000000000000010",
45331 => "0000000000000010",45332 => "0000000000000010",
45333 => "0000000000000010",45334 => "0000000000000010",
45335 => "0000000000000010",45336 => "0000000000000010",
45337 => "0000000000000010",45338 => "0000000000000010",
45339 => "0000000000000010",45340 => "0000000000000010",
45341 => "0000000000000010",45342 => "0000000000000010",
45343 => "0000000000000010",45344 => "0000000000000010",
45345 => "0000000000000010",45346 => "0000000000000010",
45347 => "0000000000000010",45348 => "0000000000000010",
45349 => "0000000000000010",45350 => "0000000000000010",
45351 => "0000000000000010",45352 => "0000000000000010",
45353 => "0000000000000010",45354 => "0000000000000010",
45355 => "0000000000000010",45356 => "0000000000000010",
45357 => "0000000000000010",45358 => "0000000000000010",
45359 => "0000000000000010",45360 => "0000000000000010",
45361 => "0000000000000010",45362 => "0000000000000010",
45363 => "0000000000000010",45364 => "0000000000000010",
45365 => "0000000000000010",45366 => "0000000000000010",
45367 => "0000000000000010",45368 => "0000000000000010",
45369 => "0000000000000010",45370 => "0000000000000010",
45371 => "0000000000000010",45372 => "0000000000000010",
45373 => "0000000000000010",45374 => "0000000000000010",
45375 => "0000000000000010",45376 => "0000000000000010",
45377 => "0000000000000010",45378 => "0000000000000010",
45379 => "0000000000000010",45380 => "0000000000000010",
45381 => "0000000000000010",45382 => "0000000000000010",
45383 => "0000000000000010",45384 => "0000000000000010",
45385 => "0000000000000010",45386 => "0000000000000010",
45387 => "0000000000000010",45388 => "0000000000000010",
45389 => "0000000000000010",45390 => "0000000000000010",
45391 => "0000000000000010",45392 => "0000000000000010",
45393 => "0000000000000010",45394 => "0000000000000010",
45395 => "0000000000000010",45396 => "0000000000000010",
45397 => "0000000000000010",45398 => "0000000000000010",
45399 => "0000000000000010",45400 => "0000000000000010",
45401 => "0000000000000010",45402 => "0000000000000010",
45403 => "0000000000000010",45404 => "0000000000000010",
45405 => "0000000000000010",45406 => "0000000000000010",
45407 => "0000000000000010",45408 => "0000000000000010",
45409 => "0000000000000010",45410 => "0000000000000010",
45411 => "0000000000000010",45412 => "0000000000000010",
45413 => "0000000000000010",45414 => "0000000000000010",
45415 => "0000000000000010",45416 => "0000000000000010",
45417 => "0000000000000010",45418 => "0000000000000010",
45419 => "0000000000000010",45420 => "0000000000000010",
45421 => "0000000000000010",45422 => "0000000000000010",
45423 => "0000000000000010",45424 => "0000000000000010",
45425 => "0000000000000010",45426 => "0000000000000010",
45427 => "0000000000000010",45428 => "0000000000000010",
45429 => "0000000000000010",45430 => "0000000000000010",
45431 => "0000000000000010",45432 => "0000000000000010",
45433 => "0000000000000010",45434 => "0000000000000010",
45435 => "0000000000000010",45436 => "0000000000000010",
45437 => "0000000000000010",45438 => "0000000000000010",
45439 => "0000000000000010",45440 => "0000000000000010",
45441 => "0000000000000010",45442 => "0000000000000010",
45443 => "0000000000000010",45444 => "0000000000000010",
45445 => "0000000000000010",45446 => "0000000000000010",
45447 => "0000000000000010",45448 => "0000000000000010",
45449 => "0000000000000010",45450 => "0000000000000010",
45451 => "0000000000000010",45452 => "0000000000000010",
45453 => "0000000000000010",45454 => "0000000000000010",
45455 => "0000000000000010",45456 => "0000000000000010",
45457 => "0000000000000010",45458 => "0000000000000010",
45459 => "0000000000000010",45460 => "0000000000000010",
45461 => "0000000000000010",45462 => "0000000000000010",
45463 => "0000000000000010",45464 => "0000000000000010",
45465 => "0000000000000010",45466 => "0000000000000010",
45467 => "0000000000000010",45468 => "0000000000000010",
45469 => "0000000000000010",45470 => "0000000000000010",
45471 => "0000000000000010",45472 => "0000000000000010",
45473 => "0000000000000010",45474 => "0000000000000010",
45475 => "0000000000000010",45476 => "0000000000000010",
45477 => "0000000000000010",45478 => "0000000000000010",
45479 => "0000000000000010",45480 => "0000000000000010",
45481 => "0000000000000010",45482 => "0000000000000010",
45483 => "0000000000000010",45484 => "0000000000000010",
45485 => "0000000000000010",45486 => "0000000000000010",
45487 => "0000000000000010",45488 => "0000000000000010",
45489 => "0000000000000010",45490 => "0000000000000010",
45491 => "0000000000000010",45492 => "0000000000000010",
45493 => "0000000000000010",45494 => "0000000000000010",
45495 => "0000000000000010",45496 => "0000000000000010",
45497 => "0000000000000010",45498 => "0000000000000010",
45499 => "0000000000000010",45500 => "0000000000000010",
45501 => "0000000000000010",45502 => "0000000000000010",
45503 => "0000000000000010",45504 => "0000000000000010",
45505 => "0000000000000010",45506 => "0000000000000010",
45507 => "0000000000000010",45508 => "0000000000000010",
45509 => "0000000000000010",45510 => "0000000000000010",
45511 => "0000000000000010",45512 => "0000000000000010",
45513 => "0000000000000010",45514 => "0000000000000010",
45515 => "0000000000000010",45516 => "0000000000000010",
45517 => "0000000000000010",45518 => "0000000000000010",
45519 => "0000000000000010",45520 => "0000000000000010",
45521 => "0000000000000010",45522 => "0000000000000010",
45523 => "0000000000000010",45524 => "0000000000000010",
45525 => "0000000000000010",45526 => "0000000000000010",
45527 => "0000000000000010",45528 => "0000000000000010",
45529 => "0000000000000010",45530 => "0000000000000010",
45531 => "0000000000000010",45532 => "0000000000000010",
45533 => "0000000000000010",45534 => "0000000000000010",
45535 => "0000000000000010",45536 => "0000000000000010",
45537 => "0000000000000010",45538 => "0000000000000010",
45539 => "0000000000000010",45540 => "0000000000000010",
45541 => "0000000000000010",45542 => "0000000000000010",
45543 => "0000000000000010",45544 => "0000000000000010",
45545 => "0000000000000010",45546 => "0000000000000010",
45547 => "0000000000000010",45548 => "0000000000000010",
45549 => "0000000000000010",45550 => "0000000000000010",
45551 => "0000000000000010",45552 => "0000000000000010",
45553 => "0000000000000010",45554 => "0000000000000010",
45555 => "0000000000000010",45556 => "0000000000000010",
45557 => "0000000000000010",45558 => "0000000000000010",
45559 => "0000000000000001",45560 => "0000000000000001",
45561 => "0000000000000001",45562 => "0000000000000001",
45563 => "0000000000000001",45564 => "0000000000000001",
45565 => "0000000000000001",45566 => "0000000000000001",
45567 => "0000000000000001",45568 => "0000000000000001",
45569 => "0000000000000001",45570 => "0000000000000001",
45571 => "0000000000000001",45572 => "0000000000000001",
45573 => "0000000000000001",45574 => "0000000000000001",
45575 => "0000000000000001",45576 => "0000000000000001",
45577 => "0000000000000001",45578 => "0000000000000001",
45579 => "0000000000000001",45580 => "0000000000000001",
45581 => "0000000000000001",45582 => "0000000000000001",
45583 => "0000000000000001",45584 => "0000000000000001",
45585 => "0000000000000001",45586 => "0000000000000001",
45587 => "0000000000000001",45588 => "0000000000000001",
45589 => "0000000000000001",45590 => "0000000000000001",
45591 => "0000000000000001",45592 => "0000000000000001",
45593 => "0000000000000001",45594 => "0000000000000001",
45595 => "0000000000000001",45596 => "0000000000000001",
45597 => "0000000000000001",45598 => "0000000000000001",
45599 => "0000000000000001",45600 => "0000000000000001",
45601 => "0000000000000001",45602 => "0000000000000001",
45603 => "0000000000000001",45604 => "0000000000000001",
45605 => "0000000000000001",45606 => "0000000000000001",
45607 => "0000000000000001",45608 => "0000000000000001",
45609 => "0000000000000001",45610 => "0000000000000001",
45611 => "0000000000000001",45612 => "0000000000000001",
45613 => "0000000000000001",45614 => "0000000000000001",
45615 => "0000000000000001",45616 => "0000000000000001",
45617 => "0000000000000001",45618 => "0000000000000001",
45619 => "0000000000000001",45620 => "0000000000000001",
45621 => "0000000000000001",45622 => "0000000000000001",
45623 => "0000000000000001",45624 => "0000000000000001",
45625 => "0000000000000001",45626 => "0000000000000001",
45627 => "0000000000000001",45628 => "0000000000000001",
45629 => "0000000000000001",45630 => "0000000000000001",
45631 => "0000000000000001",45632 => "0000000000000001",
45633 => "0000000000000001",45634 => "0000000000000001",
45635 => "0000000000000001",45636 => "0000000000000001",
45637 => "0000000000000001",45638 => "0000000000000001",
45639 => "0000000000000001",45640 => "0000000000000001",
45641 => "0000000000000001",45642 => "0000000000000001",
45643 => "0000000000000001",45644 => "0000000000000001",
45645 => "0000000000000001",45646 => "0000000000000001",
45647 => "0000000000000001",45648 => "0000000000000001",
45649 => "0000000000000001",45650 => "0000000000000001",
45651 => "0000000000000001",45652 => "0000000000000001",
45653 => "0000000000000001",45654 => "0000000000000001",
45655 => "0000000000000001",45656 => "0000000000000001",
45657 => "0000000000000001",45658 => "0000000000000001",
45659 => "0000000000000001",45660 => "0000000000000001",
45661 => "0000000000000001",45662 => "0000000000000001",
45663 => "0000000000000001",45664 => "0000000000000001",
45665 => "0000000000000001",45666 => "0000000000000001",
45667 => "0000000000000001",45668 => "0000000000000001",
45669 => "0000000000000001",45670 => "0000000000000001",
45671 => "0000000000000001",45672 => "0000000000000001",
45673 => "0000000000000001",45674 => "0000000000000001",
45675 => "0000000000000001",45676 => "0000000000000001",
45677 => "0000000000000001",45678 => "0000000000000001",
45679 => "0000000000000001",45680 => "0000000000000001",
45681 => "0000000000000001",45682 => "0000000000000001",
45683 => "0000000000000001",45684 => "0000000000000001",
45685 => "0000000000000001",45686 => "0000000000000001",
45687 => "0000000000000001",45688 => "0000000000000001",
45689 => "0000000000000001",45690 => "0000000000000001",
45691 => "0000000000000001",45692 => "0000000000000001",
45693 => "0000000000000001",45694 => "0000000000000001",
45695 => "0000000000000001",45696 => "0000000000000001",
45697 => "0000000000000001",45698 => "0000000000000001",
45699 => "0000000000000001",45700 => "0000000000000001",
45701 => "0000000000000001",45702 => "0000000000000001",
45703 => "0000000000000001",45704 => "0000000000000001",
45705 => "0000000000000001",45706 => "0000000000000001",
45707 => "0000000000000001",45708 => "0000000000000001",
45709 => "0000000000000001",45710 => "0000000000000001",
45711 => "0000000000000001",45712 => "0000000000000001",
45713 => "0000000000000001",45714 => "0000000000000001",
45715 => "0000000000000001",45716 => "0000000000000001",
45717 => "0000000000000001",45718 => "0000000000000001",
45719 => "0000000000000001",45720 => "0000000000000001",
45721 => "0000000000000001",45722 => "0000000000000001",
45723 => "0000000000000001",45724 => "0000000000000001",
45725 => "0000000000000001",45726 => "0000000000000001",
45727 => "0000000000000001",45728 => "0000000000000001",
45729 => "0000000000000001",45730 => "0000000000000001",
45731 => "0000000000000001",45732 => "0000000000000001",
45733 => "0000000000000001",45734 => "0000000000000001",
45735 => "0000000000000001",45736 => "0000000000000001",
45737 => "0000000000000001",45738 => "0000000000000001",
45739 => "0000000000000001",45740 => "0000000000000001",
45741 => "0000000000000001",45742 => "0000000000000001",
45743 => "0000000000000001",45744 => "0000000000000001",
45745 => "0000000000000001",45746 => "0000000000000001",
45747 => "0000000000000001",45748 => "0000000000000001",
45749 => "0000000000000001",45750 => "0000000000000001",
45751 => "0000000000000001",45752 => "0000000000000001",
45753 => "0000000000000001",45754 => "0000000000000001",
45755 => "0000000000000001",45756 => "0000000000000001",
45757 => "0000000000000001",45758 => "0000000000000001",
45759 => "0000000000000001",45760 => "0000000000000001",
45761 => "0000000000000001",45762 => "0000000000000001",
45763 => "0000000000000001",45764 => "0000000000000001",
45765 => "0000000000000001",45766 => "0000000000000001",
45767 => "0000000000000001",45768 => "0000000000000001",
45769 => "0000000000000001",45770 => "0000000000000001",
45771 => "0000000000000001",45772 => "0000000000000001",
45773 => "0000000000000001",45774 => "0000000000000001",
45775 => "0000000000000001",45776 => "0000000000000001",
45777 => "0000000000000001",45778 => "0000000000000001",
45779 => "0000000000000001",45780 => "0000000000000001",
45781 => "0000000000000001",45782 => "0000000000000001",
45783 => "0000000000000001",45784 => "0000000000000001",
45785 => "0000000000000001",45786 => "0000000000000001",
45787 => "0000000000000001",45788 => "0000000000000001",
45789 => "0000000000000001",45790 => "0000000000000001",
45791 => "0000000000000001",45792 => "0000000000000001",
45793 => "0000000000000001",45794 => "0000000000000001",
45795 => "0000000000000001",45796 => "0000000000000001",
45797 => "0000000000000001",45798 => "0000000000000001",
45799 => "0000000000000001",45800 => "0000000000000001",
45801 => "0000000000000001",45802 => "0000000000000001",
45803 => "0000000000000001",45804 => "0000000000000001",
45805 => "0000000000000001",45806 => "0000000000000001",
45807 => "0000000000000001",45808 => "0000000000000001",
45809 => "0000000000000001",45810 => "0000000000000001",
45811 => "0000000000000001",45812 => "0000000000000001",
45813 => "0000000000000001",45814 => "0000000000000001",
45815 => "0000000000000001",45816 => "0000000000000001",
45817 => "0000000000000001",45818 => "0000000000000001",
45819 => "0000000000000001",45820 => "0000000000000001",
45821 => "0000000000000001",45822 => "0000000000000001",
45823 => "0000000000000001",45824 => "0000000000000001",
45825 => "0000000000000001",45826 => "0000000000000001",
45827 => "0000000000000001",45828 => "0000000000000001",
45829 => "0000000000000001",45830 => "0000000000000001",
45831 => "0000000000000001",45832 => "0000000000000001",
45833 => "0000000000000001",45834 => "0000000000000001",
45835 => "0000000000000001",45836 => "0000000000000001",
45837 => "0000000000000001",45838 => "0000000000000001",
45839 => "0000000000000001",45840 => "0000000000000001",
45841 => "0000000000000001",45842 => "0000000000000001",
45843 => "0000000000000001",45844 => "0000000000000001",
45845 => "0000000000000001",45846 => "0000000000000001",
45847 => "0000000000000001",45848 => "0000000000000001",
45849 => "0000000000000001",45850 => "0000000000000001",
45851 => "0000000000000001",45852 => "0000000000000001",
45853 => "0000000000000001",45854 => "0000000000000001",
45855 => "0000000000000001",45856 => "0000000000000001",
45857 => "0000000000000001",45858 => "0000000000000001",
45859 => "0000000000000001",45860 => "0000000000000001",
45861 => "0000000000000001",45862 => "0000000000000001",
45863 => "0000000000000001",45864 => "0000000000000001",
45865 => "0000000000000001",45866 => "0000000000000001",
45867 => "0000000000000001",45868 => "0000000000000001",
45869 => "0000000000000001",45870 => "0000000000000001",
45871 => "0000000000000001",45872 => "0000000000000001",
45873 => "0000000000000001",45874 => "0000000000000001",
45875 => "0000000000000001",45876 => "0000000000000001",
45877 => "0000000000000001",45878 => "0000000000000001",
45879 => "0000000000000001",45880 => "0000000000000001",
45881 => "0000000000000001",45882 => "0000000000000001",
45883 => "0000000000000001",45884 => "0000000000000001",
45885 => "0000000000000001",45886 => "0000000000000001",
45887 => "0000000000000001",45888 => "0000000000000001",
45889 => "0000000000000001",45890 => "0000000000000001",
45891 => "0000000000000001",45892 => "0000000000000001",
45893 => "0000000000000001",45894 => "0000000000000001",
45895 => "0000000000000001",45896 => "0000000000000001",
45897 => "0000000000000001",45898 => "0000000000000001",
45899 => "0000000000000001",45900 => "0000000000000001",
45901 => "0000000000000001",45902 => "0000000000000001",
45903 => "0000000000000001",45904 => "0000000000000001",
45905 => "0000000000000001",45906 => "0000000000000001",
45907 => "0000000000000001",45908 => "0000000000000001",
45909 => "0000000000000001",45910 => "0000000000000001",
45911 => "0000000000000001",45912 => "0000000000000001",
45913 => "0000000000000001",45914 => "0000000000000001",
45915 => "0000000000000001",45916 => "0000000000000001",
45917 => "0000000000000001",45918 => "0000000000000001",
45919 => "0000000000000001",45920 => "0000000000000001",
45921 => "0000000000000001",45922 => "0000000000000001",
45923 => "0000000000000001",45924 => "0000000000000001",
45925 => "0000000000000001",45926 => "0000000000000001",
45927 => "0000000000000001",45928 => "0000000000000001",
45929 => "0000000000000001",45930 => "0000000000000001",
45931 => "0000000000000001",45932 => "0000000000000001",
45933 => "0000000000000001",45934 => "0000000000000001",
45935 => "0000000000000001",45936 => "0000000000000001",
45937 => "0000000000000001",45938 => "0000000000000001",
45939 => "0000000000000001",45940 => "0000000000000001",
45941 => "0000000000000001",45942 => "0000000000000001",
45943 => "0000000000000001",45944 => "0000000000000001",
45945 => "0000000000000001",45946 => "0000000000000001",
45947 => "0000000000000001",45948 => "0000000000000001",
45949 => "0000000000000001",45950 => "0000000000000001",
45951 => "0000000000000001",45952 => "0000000000000001",
45953 => "0000000000000001",45954 => "0000000000000001",
45955 => "0000000000000001",45956 => "0000000000000001",
45957 => "0000000000000001",45958 => "0000000000000001",
45959 => "0000000000000001",45960 => "0000000000000001",
45961 => "0000000000000001",45962 => "0000000000000001",
45963 => "0000000000000001",45964 => "0000000000000001",
45965 => "0000000000000001",45966 => "0000000000000001",
45967 => "0000000000000001",45968 => "0000000000000001",
45969 => "0000000000000001",45970 => "0000000000000001",
45971 => "0000000000000001",45972 => "0000000000000001",
45973 => "0000000000000001",45974 => "0000000000000001",
45975 => "0000000000000001",45976 => "0000000000000001",
45977 => "0000000000000001",45978 => "0000000000000001",
45979 => "0000000000000001",45980 => "0000000000000001",
45981 => "0000000000000001",45982 => "0000000000000001",
45983 => "0000000000000001",45984 => "0000000000000001",
45985 => "0000000000000001",45986 => "0000000000000001",
45987 => "0000000000000001",45988 => "0000000000000001",
45989 => "0000000000000001",45990 => "0000000000000001",
45991 => "0000000000000001",45992 => "0000000000000001",
45993 => "0000000000000001",45994 => "0000000000000001",
45995 => "0000000000000001",45996 => "0000000000000001",
45997 => "0000000000000001",45998 => "0000000000000001",
45999 => "0000000000000001",46000 => "0000000000000001",
46001 => "0000000000000001",46002 => "0000000000000001",
46003 => "0000000000000001",46004 => "0000000000000001",
46005 => "0000000000000001",46006 => "0000000000000001",
46007 => "0000000000000001",46008 => "0000000000000001",
46009 => "0000000000000001",46010 => "0000000000000001",
46011 => "0000000000000001",46012 => "0000000000000001",
46013 => "0000000000000001",46014 => "0000000000000001",
46015 => "0000000000000001",46016 => "0000000000000001",
46017 => "0000000000000001",46018 => "0000000000000001",
46019 => "0000000000000001",46020 => "0000000000000001",
46021 => "0000000000000001",46022 => "0000000000000001",
46023 => "0000000000000001",46024 => "0000000000000001",
46025 => "0000000000000001",46026 => "0000000000000001",
46027 => "0000000000000001",46028 => "0000000000000001",
46029 => "0000000000000001",46030 => "0000000000000001",
46031 => "0000000000000001",46032 => "0000000000000001",
46033 => "0000000000000001",46034 => "0000000000000001",
46035 => "0000000000000001",46036 => "0000000000000001",
46037 => "0000000000000001",46038 => "0000000000000001",
46039 => "0000000000000001",46040 => "0000000000000001",
46041 => "0000000000000001",46042 => "0000000000000001",
46043 => "0000000000000001",46044 => "0000000000000001",
46045 => "0000000000000001",46046 => "0000000000000001",
46047 => "0000000000000001",46048 => "0000000000000001",
46049 => "0000000000000001",46050 => "0000000000000001",
46051 => "0000000000000001",46052 => "0000000000000001",
46053 => "0000000000000001",46054 => "0000000000000001",
46055 => "0000000000000001",46056 => "0000000000000010",
46057 => "0000000000000010",46058 => "0000000000000010",
46059 => "0000000000000010",46060 => "0000000000000010",
46061 => "0000000000000010",46062 => "0000000000000010",
46063 => "0000000000000010",46064 => "0000000000000010",
46065 => "0000000000000010",46066 => "0000000000000010",
46067 => "0000000000000010",46068 => "0000000000000010",
46069 => "0000000000000010",46070 => "0000000000000010",
46071 => "0000000000000010",46072 => "0000000000000010",
46073 => "0000000000000010",46074 => "0000000000000010",
46075 => "0000000000000010",46076 => "0000000000000010",
46077 => "0000000000000010",46078 => "0000000000000010",
46079 => "0000000000000010",46080 => "0000000000000010",
46081 => "0000000000000010",46082 => "0000000000000010",
46083 => "0000000000000010",46084 => "0000000000000010",
46085 => "0000000000000010",46086 => "0000000000000010",
46087 => "0000000000000010",46088 => "0000000000000010",
46089 => "0000000000000010",46090 => "0000000000000010",
46091 => "0000000000000010",46092 => "0000000000000010",
46093 => "0000000000000010",46094 => "0000000000000010",
46095 => "0000000000000010",46096 => "0000000000000010",
46097 => "0000000000000010",46098 => "0000000000000010",
46099 => "0000000000000010",46100 => "0000000000000010",
46101 => "0000000000000010",46102 => "0000000000000010",
46103 => "0000000000000010",46104 => "0000000000000010",
46105 => "0000000000000010",46106 => "0000000000000010",
46107 => "0000000000000010",46108 => "0000000000000010",
46109 => "0000000000000010",46110 => "0000000000000010",
46111 => "0000000000000010",46112 => "0000000000000010",
46113 => "0000000000000010",46114 => "0000000000000010",
46115 => "0000000000000010",46116 => "0000000000000010",
46117 => "0000000000000010",46118 => "0000000000000010",
46119 => "0000000000000010",46120 => "0000000000000010",
46121 => "0000000000000010",46122 => "0000000000000010",
46123 => "0000000000000010",46124 => "0000000000000010",
46125 => "0000000000000010",46126 => "0000000000000010",
46127 => "0000000000000010",46128 => "0000000000000010",
46129 => "0000000000000010",46130 => "0000000000000010",
46131 => "0000000000000010",46132 => "0000000000000010",
46133 => "0000000000000010",46134 => "0000000000000010",
46135 => "0000000000000010",46136 => "0000000000000010",
46137 => "0000000000000010",46138 => "0000000000000010",
46139 => "0000000000000010",46140 => "0000000000000010",
46141 => "0000000000000010",46142 => "0000000000000010",
46143 => "0000000000000010",46144 => "0000000000000010",
46145 => "0000000000000010",46146 => "0000000000000010",
46147 => "0000000000000010",46148 => "0000000000000010",
46149 => "0000000000000010",46150 => "0000000000000010",
46151 => "0000000000000010",46152 => "0000000000000010",
46153 => "0000000000000010",46154 => "0000000000000010",
46155 => "0000000000000010",46156 => "0000000000000010",
46157 => "0000000000000010",46158 => "0000000000000010",
46159 => "0000000000000010",46160 => "0000000000000010",
46161 => "0000000000000010",46162 => "0000000000000010",
46163 => "0000000000000010",46164 => "0000000000000010",
46165 => "0000000000000010",46166 => "0000000000000010",
46167 => "0000000000000010",46168 => "0000000000000010",
46169 => "0000000000000010",46170 => "0000000000000010",
46171 => "0000000000000010",46172 => "0000000000000010",
46173 => "0000000000000010",46174 => "0000000000000010",
46175 => "0000000000000010",46176 => "0000000000000010",
46177 => "0000000000000010",46178 => "0000000000000010",
46179 => "0000000000000010",46180 => "0000000000000010",
46181 => "0000000000000010",46182 => "0000000000000010",
46183 => "0000000000000010",46184 => "0000000000000010",
46185 => "0000000000000010",46186 => "0000000000000010",
46187 => "0000000000000010",46188 => "0000000000000010",
46189 => "0000000000000010",46190 => "0000000000000010",
46191 => "0000000000000010",46192 => "0000000000000010",
46193 => "0000000000000010",46194 => "0000000000000010",
46195 => "0000000000000010",46196 => "0000000000000010",
46197 => "0000000000000010",46198 => "0000000000000010",
46199 => "0000000000000010",46200 => "0000000000000010",
46201 => "0000000000000010",46202 => "0000000000000010",
46203 => "0000000000000010",46204 => "0000000000000010",
46205 => "0000000000000010",46206 => "0000000000000010",
46207 => "0000000000000010",46208 => "0000000000000010",
46209 => "0000000000000010",46210 => "0000000000000010",
46211 => "0000000000000010",46212 => "0000000000000010",
46213 => "0000000000000010",46214 => "0000000000000010",
46215 => "0000000000000010",46216 => "0000000000000010",
46217 => "0000000000000010",46218 => "0000000000000010",
46219 => "0000000000000010",46220 => "0000000000000010",
46221 => "0000000000000010",46222 => "0000000000000010",
46223 => "0000000000000010",46224 => "0000000000000010",
46225 => "0000000000000010",46226 => "0000000000000010",
46227 => "0000000000000010",46228 => "0000000000000010",
46229 => "0000000000000010",46230 => "0000000000000010",
46231 => "0000000000000010",46232 => "0000000000000010",
46233 => "0000000000000010",46234 => "0000000000000010",
46235 => "0000000000000010",46236 => "0000000000000010",
46237 => "0000000000000010",46238 => "0000000000000010",
46239 => "0000000000000010",46240 => "0000000000000010",
46241 => "0000000000000010",46242 => "0000000000000010",
46243 => "0000000000000010",46244 => "0000000000000010",
46245 => "0000000000000010",46246 => "0000000000000010",
46247 => "0000000000000010",46248 => "0000000000000010",
46249 => "0000000000000010",46250 => "0000000000000010",
46251 => "0000000000000010",46252 => "0000000000000010",
46253 => "0000000000000010",46254 => "0000000000000010",
46255 => "0000000000000010",46256 => "0000000000000010",
46257 => "0000000000000010",46258 => "0000000000000010",
46259 => "0000000000000010",46260 => "0000000000000010",
46261 => "0000000000000010",46262 => "0000000000000010",
46263 => "0000000000000010",46264 => "0000000000000010",
46265 => "0000000000000010",46266 => "0000000000000010",
46267 => "0000000000000010",46268 => "0000000000000010",
46269 => "0000000000000010",46270 => "0000000000000010",
46271 => "0000000000000010",46272 => "0000000000000010",
46273 => "0000000000000010",46274 => "0000000000000010",
46275 => "0000000000000010",46276 => "0000000000000010",
46277 => "0000000000000010",46278 => "0000000000000010",
46279 => "0000000000000010",46280 => "0000000000000010",
46281 => "0000000000000010",46282 => "0000000000000010",
46283 => "0000000000000010",46284 => "0000000000000010",
46285 => "0000000000000010",46286 => "0000000000000010",
46287 => "0000000000000010",46288 => "0000000000000010",
46289 => "0000000000000010",46290 => "0000000000000010",
46291 => "0000000000000010",46292 => "0000000000000010",
46293 => "0000000000000010",46294 => "0000000000000010",
46295 => "0000000000000010",46296 => "0000000000000010",
46297 => "0000000000000010",46298 => "0000000000000010",
46299 => "0000000000000010",46300 => "0000000000000010",
46301 => "0000000000000010",46302 => "0000000000000010",
46303 => "0000000000000010",46304 => "0000000000000010",
46305 => "0000000000000010",46306 => "0000000000000010",
46307 => "0000000000000010",46308 => "0000000000000010",
46309 => "0000000000000010",46310 => "0000000000000010",
46311 => "0000000000000010",46312 => "0000000000000010",
46313 => "0000000000000010",46314 => "0000000000000010",
46315 => "0000000000000010",46316 => "0000000000000010",
46317 => "0000000000000010",46318 => "0000000000000010",
46319 => "0000000000000010",46320 => "0000000000000010",
46321 => "0000000000000010",46322 => "0000000000000010",
46323 => "0000000000000010",46324 => "0000000000000010",
46325 => "0000000000000010",46326 => "0000000000000010",
46327 => "0000000000000010",46328 => "0000000000000010",
46329 => "0000000000000010",46330 => "0000000000000010",
46331 => "0000000000000010",46332 => "0000000000000010",
46333 => "0000000000000010",46334 => "0000000000000010",
46335 => "0000000000000010",46336 => "0000000000000010",
46337 => "0000000000000010",46338 => "0000000000000010",
46339 => "0000000000000010",46340 => "0000000000000010",
46341 => "0000000000000010",46342 => "0000000000000010",
46343 => "0000000000000010",46344 => "0000000000000010",
46345 => "0000000000000010",46346 => "0000000000000010",
46347 => "0000000000000010",46348 => "0000000000000010",
46349 => "0000000000000010",46350 => "0000000000000010",
46351 => "0000000000000010",46352 => "0000000000000010",
46353 => "0000000000000010",46354 => "0000000000000010",
46355 => "0000000000000010",46356 => "0000000000000010",
46357 => "0000000000000010",46358 => "0000000000000010",
46359 => "0000000000000010",46360 => "0000000000000010",
46361 => "0000000000000010",46362 => "0000000000000010",
46363 => "0000000000000010",46364 => "0000000000000010",
46365 => "0000000000000010",46366 => "0000000000000010",
46367 => "0000000000000010",46368 => "0000000000000010",
46369 => "0000000000000010",46370 => "0000000000000010",
46371 => "0000000000000010",46372 => "0000000000000010",
46373 => "0000000000000010",46374 => "0000000000000010",
46375 => "0000000000000010",46376 => "0000000000000010",
46377 => "0000000000000010",46378 => "0000000000000010",
46379 => "0000000000000010",46380 => "0000000000000010",
46381 => "0000000000000010",46382 => "0000000000000010",
46383 => "0000000000000010",46384 => "0000000000000010",
46385 => "0000000000000010",46386 => "0000000000000010",
46387 => "0000000000000010",46388 => "0000000000000010",
46389 => "0000000000000010",46390 => "0000000000000010",
46391 => "0000000000000010",46392 => "0000000000000010",
46393 => "0000000000000010",46394 => "0000000000000010",
46395 => "0000000000000010",46396 => "0000000000000010",
46397 => "0000000000000010",46398 => "0000000000000010",
46399 => "0000000000000010",46400 => "0000000000000010",
46401 => "0000000000000010",46402 => "0000000000000010",
46403 => "0000000000000010",46404 => "0000000000000010",
46405 => "0000000000000010",46406 => "0000000000000010",
46407 => "0000000000000010",46408 => "0000000000000010",
46409 => "0000000000000010",46410 => "0000000000000010",
46411 => "0000000000000010",46412 => "0000000000000010",
46413 => "0000000000000010",46414 => "0000000000000010",
46415 => "0000000000000010",46416 => "0000000000000010",
46417 => "0000000000000010",46418 => "0000000000000010",
46419 => "0000000000000010",46420 => "0000000000000010",
46421 => "0000000000000010",46422 => "0000000000000010",
46423 => "0000000000000010",46424 => "0000000000000010",
46425 => "0000000000000010",46426 => "0000000000000010",
46427 => "0000000000000010",46428 => "0000000000000010",
46429 => "0000000000000010",46430 => "0000000000000010",
46431 => "0000000000000010",46432 => "0000000000000010",
46433 => "0000000000000010",46434 => "0000000000000010",
46435 => "0000000000000010",46436 => "0000000000000010",
46437 => "0000000000000010",46438 => "0000000000000010",
46439 => "0000000000000010",46440 => "0000000000000010",
46441 => "0000000000000010",46442 => "0000000000000010",
46443 => "0000000000000010",46444 => "0000000000000010",
46445 => "0000000000000010",46446 => "0000000000000010",
46447 => "0000000000000010",46448 => "0000000000000010",
46449 => "0000000000000010",46450 => "0000000000000010",
46451 => "0000000000000010",46452 => "0000000000000010",
46453 => "0000000000000010",46454 => "0000000000000010",
46455 => "0000000000000010",46456 => "0000000000000010",
46457 => "0000000000000010",46458 => "0000000000000010",
46459 => "0000000000000010",46460 => "0000000000000010",
46461 => "0000000000000010",46462 => "0000000000000010",
46463 => "0000000000000010",46464 => "0000000000000010",
46465 => "0000000000000010",46466 => "0000000000000010",
46467 => "0000000000000010",46468 => "0000000000000010",
46469 => "0000000000000010",46470 => "0000000000000010",
46471 => "0000000000000010",46472 => "0000000000000010",
46473 => "0000000000000010",46474 => "0000000000000010",
46475 => "0000000000000010",46476 => "0000000000000010",
46477 => "0000000000000010",46478 => "0000000000000010",
46479 => "0000000000000010",46480 => "0000000000000010",
46481 => "0000000000000010",46482 => "0000000000000010",
46483 => "0000000000000010",46484 => "0000000000000010",
46485 => "0000000000000010",46486 => "0000000000000010",
46487 => "0000000000000010",46488 => "0000000000000010",
46489 => "0000000000000010",46490 => "0000000000000010",
46491 => "0000000000000010",46492 => "0000000000000010",
46493 => "0000000000000010",46494 => "0000000000000010",
46495 => "0000000000000010",46496 => "0000000000000010",
46497 => "0000000000000010",46498 => "0000000000000010",
46499 => "0000000000000010",46500 => "0000000000000010",
46501 => "0000000000000010",46502 => "0000000000000010",
46503 => "0000000000000010",46504 => "0000000000000010",
46505 => "0000000000000010",46506 => "0000000000000010",
46507 => "0000000000000010",46508 => "0000000000000010",
46509 => "0000000000000010",46510 => "0000000000000010",
46511 => "0000000000000010",46512 => "0000000000000010",
46513 => "0000000000000010",46514 => "0000000000000010",
46515 => "0000000000000010",46516 => "0000000000000010",
46517 => "0000000000000010",46518 => "0000000000000010",
46519 => "0000000000000010",46520 => "0000000000000010",
46521 => "0000000000000010",46522 => "0000000000000010",
46523 => "0000000000000010",46524 => "0000000000000010",
46525 => "0000000000000010",46526 => "0000000000000010",
46527 => "0000000000000010",46528 => "0000000000000010",
46529 => "0000000000000010",46530 => "0000000000000010",
46531 => "0000000000000010",46532 => "0000000000000010",
46533 => "0000000000000010",46534 => "0000000000000010",
46535 => "0000000000000010",46536 => "0000000000000010",
46537 => "0000000000000010",46538 => "0000000000000010",
46539 => "0000000000000010",46540 => "0000000000000010",
46541 => "0000000000000010",46542 => "0000000000000010",
46543 => "0000000000000010",46544 => "0000000000000010",
46545 => "0000000000000010",46546 => "0000000000000010",
46547 => "0000000000000010",46548 => "0000000000000010",
46549 => "0000000000000010",46550 => "0000000000000010",
46551 => "0000000000000010",46552 => "0000000000000010",
46553 => "0000000000000010",46554 => "0000000000000010",
46555 => "0000000000000010",46556 => "0000000000000010",
46557 => "0000000000000010",46558 => "0000000000000010",
46559 => "0000000000000010",46560 => "0000000000000010",
46561 => "0000000000000010",46562 => "0000000000000010",
46563 => "0000000000000010",46564 => "0000000000000010",
46565 => "0000000000000010",46566 => "0000000000000010",
46567 => "0000000000000010",46568 => "0000000000000010",
46569 => "0000000000000010",46570 => "0000000000000010",
46571 => "0000000000000010",46572 => "0000000000000010",
46573 => "0000000000000010",46574 => "0000000000000010",
46575 => "0000000000000010",46576 => "0000000000000010",
46577 => "0000000000000010",46578 => "0000000000000010",
46579 => "0000000000000010",46580 => "0000000000000010",
46581 => "0000000000000010",46582 => "0000000000000010",
46583 => "0000000000000010",46584 => "0000000000000010",
46585 => "0000000000000010",46586 => "0000000000000010",
46587 => "0000000000000010",46588 => "0000000000000010",
46589 => "0000000000000010",46590 => "0000000000000010",
46591 => "0000000000000010",46592 => "0000000000000010",
46593 => "0000000000000010",46594 => "0000000000000010",
46595 => "0000000000000010",46596 => "0000000000000010",
46597 => "0000000000000010",46598 => "0000000000000010",
46599 => "0000000000000010",46600 => "0000000000000010",
46601 => "0000000000000010",46602 => "0000000000000010",
46603 => "0000000000000010",46604 => "0000000000000010",
46605 => "0000000000000010",46606 => "0000000000000010",
46607 => "0000000000000010",46608 => "0000000000000010",
46609 => "0000000000000010",46610 => "0000000000000010",
46611 => "0000000000000010",46612 => "0000000000000010",
46613 => "0000000000000010",46614 => "0000000000000010",
46615 => "0000000000000010",46616 => "0000000000000010",
46617 => "0000000000000010",46618 => "0000000000000010",
46619 => "0000000000000010",46620 => "0000000000000010",
46621 => "0000000000000010",46622 => "0000000000000010",
46623 => "0000000000000010",46624 => "0000000000000010",
46625 => "0000000000000010",46626 => "0000000000000010",
46627 => "0000000000000010",46628 => "0000000000000010",
46629 => "0000000000000010",46630 => "0000000000000010",
46631 => "0000000000000010",46632 => "0000000000000010",
46633 => "0000000000000010",46634 => "0000000000000010",
46635 => "0000000000000010",46636 => "0000000000000010",
46637 => "0000000000000010",46638 => "0000000000000010",
46639 => "0000000000000010",46640 => "0000000000000010",
46641 => "0000000000000010",46642 => "0000000000000010",
46643 => "0000000000000010",46644 => "0000000000000010",
46645 => "0000000000000010",46646 => "0000000000000010",
46647 => "0000000000000010",46648 => "0000000000000010",
46649 => "0000000000000010",46650 => "0000000000000010",
46651 => "0000000000000010",46652 => "0000000000000010",
46653 => "0000000000000010",46654 => "0000000000000010",
46655 => "0000000000000010",46656 => "0000000000000010",
46657 => "0000000000000010",46658 => "0000000000000010",
46659 => "0000000000000010",46660 => "0000000000000010",
46661 => "0000000000000010",46662 => "0000000000000010",
46663 => "0000000000000010",46664 => "0000000000000010",
46665 => "0000000000000010",46666 => "0000000000000010",
46667 => "0000000000000010",46668 => "0000000000000010",
46669 => "0000000000000010",46670 => "0000000000000010",
46671 => "0000000000000010",46672 => "0000000000000010",
46673 => "0000000000000010",46674 => "0000000000000010",
46675 => "0000000000000010",46676 => "0000000000000010",
46677 => "0000000000000010",46678 => "0000000000000010",
46679 => "0000000000000010",46680 => "0000000000000010",
46681 => "0000000000000010",46682 => "0000000000000010",
46683 => "0000000000000010",46684 => "0000000000000010",
46685 => "0000000000000010",46686 => "0000000000000010",
46687 => "0000000000000010",46688 => "0000000000000010",
46689 => "0000000000000010",46690 => "0000000000000010",
46691 => "0000000000000010",46692 => "0000000000000010",
46693 => "0000000000000010",46694 => "0000000000000010",
46695 => "0000000000000010",46696 => "0000000000000010",
46697 => "0000000000000010",46698 => "0000000000000010",
46699 => "0000000000000010",46700 => "0000000000000010",
46701 => "0000000000000010",46702 => "0000000000000010",
46703 => "0000000000000010",46704 => "0000000000000010",
46705 => "0000000000000010",46706 => "0000000000000010",
46707 => "0000000000000010",46708 => "0000000000000010",
46709 => "0000000000000010",46710 => "0000000000000010",
46711 => "0000000000000010",46712 => "0000000000000010",
46713 => "0000000000000010",46714 => "0000000000000010",
46715 => "0000000000000010",46716 => "0000000000000010",
46717 => "0000000000000010",46718 => "0000000000000010",
46719 => "0000000000000010",46720 => "0000000000000010",
46721 => "0000000000000010",46722 => "0000000000000010",
46723 => "0000000000000010",46724 => "0000000000000010",
46725 => "0000000000000010",46726 => "0000000000000010",
46727 => "0000000000000010",46728 => "0000000000000010",
46729 => "0000000000000010",46730 => "0000000000000010",
46731 => "0000000000000010",46732 => "0000000000000010",
46733 => "0000000000000010",46734 => "0000000000000010",
46735 => "0000000000000010",46736 => "0000000000000010",
46737 => "0000000000000010",46738 => "0000000000000010",
46739 => "0000000000000010",46740 => "0000000000000010",
46741 => "0000000000000010",46742 => "0000000000000010",
46743 => "0000000000000010",46744 => "0000000000000010",
46745 => "0000000000000010",46746 => "0000000000000010",
46747 => "0000000000000010",46748 => "0000000000000010",
46749 => "0000000000000010",46750 => "0000000000000010",
46751 => "0000000000000010",46752 => "0000000000000010",
46753 => "0000000000000010",46754 => "0000000000000010",
46755 => "0000000000000010",46756 => "0000000000000010",
46757 => "0000000000000010",46758 => "0000000000000010",
46759 => "0000000000000010",46760 => "0000000000000010",
46761 => "0000000000000010",46762 => "0000000000000010",
46763 => "0000000000000010",46764 => "0000000000000010",
46765 => "0000000000000010",46766 => "0000000000000010",
46767 => "0000000000000010",46768 => "0000000000000010",
46769 => "0000000000000010",46770 => "0000000000000010",
46771 => "0000000000000010",46772 => "0000000000000010",
46773 => "0000000000000010",46774 => "0000000000000010",
46775 => "0000000000000010",46776 => "0000000000000010",
46777 => "0000000000000010",46778 => "0000000000000010",
46779 => "0000000000000010",46780 => "0000000000000010",
46781 => "0000000000000010",46782 => "0000000000000010",
46783 => "0000000000000010",46784 => "0000000000000010",
46785 => "0000000000000010",46786 => "0000000000000010",
46787 => "0000000000000010",46788 => "0000000000000010",
46789 => "0000000000000010",46790 => "0000000000000010",
46791 => "0000000000000010",46792 => "0000000000000010",
46793 => "0000000000000010",46794 => "0000000000000010",
46795 => "0000000000000010",46796 => "0000000000000010",
46797 => "0000000000000010",46798 => "0000000000000010",
46799 => "0000000000000010",46800 => "0000000000000010",
46801 => "0000000000000010",46802 => "0000000000000010",
46803 => "0000000000000010",46804 => "0000000000000010",
46805 => "0000000000000010",46806 => "0000000000000010",
46807 => "0000000000000010",46808 => "0000000000000010",
46809 => "0000000000000010",46810 => "0000000000000010",
46811 => "0000000000000010",46812 => "0000000000000010",
46813 => "0000000000000010",46814 => "0000000000000010",
46815 => "0000000000000010",46816 => "0000000000000010",
46817 => "0000000000000010",46818 => "0000000000000010",
46819 => "0000000000000010",46820 => "0000000000000010",
46821 => "0000000000000010",46822 => "0000000000000010",
46823 => "0000000000000010",46824 => "0000000000000010",
46825 => "0000000000000010",46826 => "0000000000000010",
46827 => "0000000000000010",46828 => "0000000000000010",
46829 => "0000000000000010",46830 => "0000000000000010",
46831 => "0000000000000010",46832 => "0000000000000010",
46833 => "0000000000000010",46834 => "0000000000000010",
46835 => "0000000000000010",46836 => "0000000000000010",
46837 => "0000000000000010",46838 => "0000000000000010",
46839 => "0000000000000010",46840 => "0000000000000010",
46841 => "0000000000000010",46842 => "0000000000000010",
46843 => "0000000000000010",46844 => "0000000000000010",
46845 => "0000000000000010",46846 => "0000000000000010",
46847 => "0000000000000010",46848 => "0000000000000010",
46849 => "0000000000000010",46850 => "0000000000000010",
46851 => "0000000000000010",46852 => "0000000000000010",
46853 => "0000000000000010",46854 => "0000000000000010",
46855 => "0000000000000010",46856 => "0000000000000010",
46857 => "0000000000000010",46858 => "0000000000000010",
46859 => "0000000000000010",46860 => "0000000000000010",
46861 => "0000000000000010",46862 => "0000000000000010",
46863 => "0000000000000010",46864 => "0000000000000010",
46865 => "0000000000000010",46866 => "0000000000000010",
46867 => "0000000000000010",46868 => "0000000000000010",
46869 => "0000000000000010",46870 => "0000000000000010",
46871 => "0000000000000010",46872 => "0000000000000010",
46873 => "0000000000000010",46874 => "0000000000000010",
46875 => "0000000000000010",46876 => "0000000000000010",
46877 => "0000000000000010",46878 => "0000000000000010",
46879 => "0000000000000010",46880 => "0000000000000010",
46881 => "0000000000000010",46882 => "0000000000000010",
46883 => "0000000000000010",46884 => "0000000000000010",
46885 => "0000000000000010",46886 => "0000000000000010",
46887 => "0000000000000010",46888 => "0000000000000010",
46889 => "0000000000000010",46890 => "0000000000000010",
46891 => "0000000000000010",46892 => "0000000000000010",
46893 => "0000000000000010",46894 => "0000000000000010",
46895 => "0000000000000010",46896 => "0000000000000010",
46897 => "0000000000000010",46898 => "0000000000000010",
46899 => "0000000000000010",46900 => "0000000000000010",
46901 => "0000000000000010",46902 => "0000000000000010",
46903 => "0000000000000010",46904 => "0000000000000010",
46905 => "0000000000000010",46906 => "0000000000000010",
46907 => "0000000000000010",46908 => "0000000000000010",
46909 => "0000000000000010",46910 => "0000000000000010",
46911 => "0000000000000010",46912 => "0000000000000010",
46913 => "0000000000000010",46914 => "0000000000000010",
46915 => "0000000000000010",46916 => "0000000000000010",
46917 => "0000000000000010",46918 => "0000000000000010",
46919 => "0000000000000010",46920 => "0000000000000010",
46921 => "0000000000000010",46922 => "0000000000000010",
46923 => "0000000000000010",46924 => "0000000000000010",
46925 => "0000000000000010",46926 => "0000000000000010",
46927 => "0000000000000010",46928 => "0000000000000010",
46929 => "0000000000000010",46930 => "0000000000000010",
46931 => "0000000000000010",46932 => "0000000000000010",
46933 => "0000000000000010",46934 => "0000000000000010",
46935 => "0000000000000010",46936 => "0000000000000010",
46937 => "0000000000000010",46938 => "0000000000000010",
46939 => "0000000000000010",46940 => "0000000000000010",
46941 => "0000000000000010",46942 => "0000000000000010",
46943 => "0000000000000010",46944 => "0000000000000010",
46945 => "0000000000000010",46946 => "0000000000000010",
46947 => "0000000000000010",46948 => "0000000000000010",
46949 => "0000000000000010",46950 => "0000000000000010",
46951 => "0000000000000010",46952 => "0000000000000010",
46953 => "0000000000000010",46954 => "0000000000000010",
46955 => "0000000000000010",46956 => "0000000000000010",
46957 => "0000000000000010",46958 => "0000000000000010",
46959 => "0000000000000010",46960 => "0000000000000010",
46961 => "0000000000000010",46962 => "0000000000000010",
46963 => "0000000000000010",46964 => "0000000000000010",
46965 => "0000000000000010",46966 => "0000000000000010",
46967 => "0000000000000010",46968 => "0000000000000010",
46969 => "0000000000000010",46970 => "0000000000000010",
46971 => "0000000000000010",46972 => "0000000000000010",
46973 => "0000000000000010",46974 => "0000000000000010",
46975 => "0000000000000010",46976 => "0000000000000010",
46977 => "0000000000000010",46978 => "0000000000000010",
46979 => "0000000000000010",46980 => "0000000000000010",
46981 => "0000000000000010",46982 => "0000000000000010",
46983 => "0000000000000010",46984 => "0000000000000010",
46985 => "0000000000000010",46986 => "0000000000000010",
46987 => "0000000000000010",46988 => "0000000000000010",
46989 => "0000000000000010",46990 => "0000000000000010",
46991 => "0000000000000010",46992 => "0000000000000010",
46993 => "0000000000000010",46994 => "0000000000000010",
46995 => "0000000000000010",46996 => "0000000000000010",
46997 => "0000000000000010",46998 => "0000000000000010",
46999 => "0000000000000010",47000 => "0000000000000010",
47001 => "0000000000000010",47002 => "0000000000000010",
47003 => "0000000000000010",47004 => "0000000000000010",
47005 => "0000000000000010",47006 => "0000000000000010",
47007 => "0000000000000010",47008 => "0000000000000010",
47009 => "0000000000000010",47010 => "0000000000000010",
47011 => "0000000000000010",47012 => "0000000000000010",
47013 => "0000000000000010",47014 => "0000000000000010",
47015 => "0000000000000010",47016 => "0000000000000010",
47017 => "0000000000000010",47018 => "0000000000000010",
47019 => "0000000000000010",47020 => "0000000000000010",
47021 => "0000000000000010",47022 => "0000000000000010",
47023 => "0000000000000010",47024 => "0000000000000010",
47025 => "0000000000000010",47026 => "0000000000000010",
47027 => "0000000000000010",47028 => "0000000000000010",
47029 => "0000000000000010",47030 => "0000000000000010",
47031 => "0000000000000010",47032 => "0000000000000010",
47033 => "0000000000000010",47034 => "0000000000000010",
47035 => "0000000000000010",47036 => "0000000000000010",
47037 => "0000000000000010",47038 => "0000000000000010",
47039 => "0000000000000010",47040 => "0000000000000010",
47041 => "0000000000000010",47042 => "0000000000000010",
47043 => "0000000000000010",47044 => "0000000000000010",
47045 => "0000000000000010",47046 => "0000000000000010",
47047 => "0000000000000010",47048 => "0000000000000010",
47049 => "0000000000000010",47050 => "0000000000000010",
47051 => "0000000000000010",47052 => "0000000000000010",
47053 => "0000000000000010",47054 => "0000000000000010",
47055 => "0000000000000010",47056 => "0000000000000010",
47057 => "0000000000000010",47058 => "0000000000000010",
47059 => "0000000000000010",47060 => "0000000000000010",
47061 => "0000000000000010",47062 => "0000000000000010",
47063 => "0000000000000010",47064 => "0000000000000010",
47065 => "0000000000000010",47066 => "0000000000000010",
47067 => "0000000000000010",47068 => "0000000000000010",
47069 => "0000000000000010",47070 => "0000000000000010",
47071 => "0000000000000010",47072 => "0000000000000010",
47073 => "0000000000000010",47074 => "0000000000000010",
47075 => "0000000000000010",47076 => "0000000000000010",
47077 => "0000000000000010",47078 => "0000000000000010",
47079 => "0000000000000010",47080 => "0000000000000010",
47081 => "0000000000000010",47082 => "0000000000000010",
47083 => "0000000000000010",47084 => "0000000000000010",
47085 => "0000000000000010",47086 => "0000000000000010",
47087 => "0000000000000010",47088 => "0000000000000010",
47089 => "0000000000000010",47090 => "0000000000000010",
47091 => "0000000000000010",47092 => "0000000000000010",
47093 => "0000000000000010",47094 => "0000000000000010",
47095 => "0000000000000010",47096 => "0000000000000010",
47097 => "0000000000000010",47098 => "0000000000000010",
47099 => "0000000000000010",47100 => "0000000000000010",
47101 => "0000000000000010",47102 => "0000000000000010",
47103 => "0000000000000010",47104 => "0000000000000001",
47105 => "0000000000000001",47106 => "0000000000000001",
47107 => "0000000000000001",47108 => "0000000000000001",
47109 => "0000000000000001",47110 => "0000000000000001",
47111 => "0000000000000000",47112 => "0000000000000000",
47113 => "0000000000000000",47114 => "0000000000000001",
47115 => "0000000000000001",47116 => "0000000000000001",
47117 => "0000000000000001",47118 => "0000000000000001",
47119 => "0000000000000001",47120 => "0000000000000001",
47121 => "0000000000000001",47122 => "0000000000000001",
47123 => "0000000000000001",47124 => "0000000000000001",
47125 => "0000000000000001",47126 => "0000000000000001",
47127 => "0000000000000001",47128 => "0000000000000001",
47129 => "0000000000000001",47130 => "0000000000000001",
47131 => "0000000000000001",47132 => "0000000000000001",
47133 => "0000000000000001",47134 => "0000000000000001",
47135 => "0000000000000001",47136 => "0000000000000001",
47137 => "0000000000000001",47138 => "0000000000000001",
47139 => "0000000000000001",47140 => "0000000000000001",
47141 => "0000000000000001",47142 => "0000000000000001",
47143 => "0000000000000001",47144 => "0000000000000001",
47145 => "0000000000000001",47146 => "0000000000000001",
47147 => "0000000000000001",47148 => "0000000000000001",
47149 => "0000000000000001",47150 => "0000000000000001",
47151 => "0000000000000001",47152 => "0000000000000001",
47153 => "0000000000000001",47154 => "0000000000000001",
47155 => "0000000000000001",47156 => "0000000000000001",
47157 => "0000000000000001",47158 => "0000000000000001",
47159 => "0000000000000001",47160 => "0000000000000001",
47161 => "0000000000000001",47162 => "0000000000000001",
47163 => "0000000000000001",47164 => "0000000000000001",
47165 => "0000000000000000",47166 => "0000000000000000",
47167 => "0000000000000000",47168 => "0000000000000000",
47169 => "0000000000000000",47170 => "0000000000000000",
47171 => "0000000000000000",47172 => "0000000000000000",
47173 => "0000000000000000",47174 => "0000000000000000",
47175 => "0000000000000000",47176 => "0000000000000000",
47177 => "0000000000000000",47178 => "0000000000000000",
47179 => "0000000000000000",47180 => "0000000000000000",
47181 => "0000000000000000",47182 => "0000000000000000",
47183 => "0000000000000000",47184 => "0000000000000000",
47185 => "0000000000000000",47186 => "0000000000000000",
47187 => "0000000000000000",47188 => "0000000000000000",
47189 => "0000000000000000",47190 => "0000000000000000",
47191 => "0000000000000000",47192 => "0000000000000000",
47193 => "0000000000000000",47194 => "0000000000000000",
47195 => "0000000000000000",47196 => "0000000000000000",
47197 => "0000000000000000",47198 => "0000000000000000",
47199 => "0000000000000000",47200 => "0000000000000000",
47201 => "0000000000000000",47202 => "0000000000000000",
47203 => "0000000000000000",47204 => "0000000000000001",
47205 => "0000000000000001",47206 => "0000000000000001",
47207 => "0000000000000001",47208 => "0000000000000001",
47209 => "0000000000000001",47210 => "0000000000000001",
47211 => "0000000000000001",47212 => "0000000000000001",
47213 => "0000000000000001",47214 => "0000000000000001",
47215 => "0000000000000001",47216 => "0000000000000001",
47217 => "0000000000000001",47218 => "0000000000000001",
47219 => "0000000000000001",47220 => "0000000000000001",
47221 => "0000000000000001",47222 => "0000000000000001",
47223 => "0000000000000001",47224 => "0000000000000001",
47225 => "0000000000000001",47226 => "0000000000000001",
47227 => "0000000000000001",47228 => "0000000000000001",
47229 => "0000000000000001",47230 => "0000000000000001",
47231 => "0000000000000001",47232 => "0000000000000001",
47233 => "0000000000000001",47234 => "0000000000000001",
47235 => "0000000000000001",47236 => "0000000000000001",
47237 => "0000000000000001",47238 => "0000000000000001",
47239 => "0000000000000001",47240 => "0000000000000001",
47241 => "0000000000000001",47242 => "0000000000000001",
47243 => "0000000000000001",47244 => "0000000000000001",
47245 => "0000000000000001",47246 => "0000000000000001",
47247 => "0000000000000001",47248 => "0000000000000001",
47249 => "0000000000000001",47250 => "0000000000000001",
47251 => "0000000000000001",47252 => "0000000000000001",
47253 => "0000000000000001",47254 => "0000000000000001",
47255 => "0000000000000001",47256 => "0000000000000001",
47257 => "0000000000000001",47258 => "0000000000000001",
47259 => "0000000000000001",47260 => "0000000000000001",
47261 => "0000000000000001",47262 => "0000000000000001",
47263 => "0000000000000001",47264 => "0000000000000001",
47265 => "0000000000000001",47266 => "0000000000000001",
47267 => "0000000000000001",47268 => "0000000000000001",
47269 => "0000000000000001",47270 => "0000000000000001",
47271 => "0000000000000001",47272 => "0000000000000001",
47273 => "0000000000000001",47274 => "0000000000000001",
47275 => "0000000000000001",47276 => "0000000000000001",
47277 => "0000000000000001",47278 => "0000000000000001",
47279 => "0000000000000001",47280 => "0000000000000001",
47281 => "0000000000000001",47282 => "0000000000000001",
47283 => "0000000000000001",47284 => "0000000000000001",
47285 => "0000000000000001",47286 => "0000000000000001",
47287 => "0000000000000001",47288 => "0000000000000001",
47289 => "0000000000000001",47290 => "0000000000000001",
47291 => "0000000000000001",47292 => "0000000000000001",
47293 => "0000000000000001",47294 => "0000000000000001",
47295 => "0000000000000001",47296 => "0000000000000001",
47297 => "0000000000000001",47298 => "0000000000000001",
47299 => "0000000000000001",47300 => "0000000000000001",
47301 => "0000000000000001",47302 => "0000000000000001",
47303 => "0000000000000001",47304 => "0000000000000001",
47305 => "0000000000000001",47306 => "0000000000000001",
47307 => "0000000000000001",47308 => "0000000000000001",
47309 => "0000000000000001",47310 => "0000000000000001",
47311 => "0000000000000001",47312 => "0000000000000001",
47313 => "0000000000000001",47314 => "0000000000000001",
47315 => "0000000000000001",47316 => "0000000000000001",
47317 => "0000000000000001",47318 => "0000000000000001",
47319 => "0000000000000001",47320 => "0000000000000001",
47321 => "0000000000000001",47322 => "0000000000000001",
47323 => "0000000000000001",47324 => "0000000000000001",
47325 => "0000000000000001",47326 => "0000000000000001",
47327 => "0000000000000001",47328 => "0000000000000001",
47329 => "0000000000000001",47330 => "0000000000000001",
47331 => "0000000000000001",47332 => "0000000000000001",
47333 => "0000000000000001",47334 => "0000000000000001",
47335 => "0000000000000001",47336 => "0000000000000001",
47337 => "0000000000000001",47338 => "0000000000000001",
47339 => "0000000000000001",47340 => "0000000000000001",
47341 => "0000000000000001",47342 => "0000000000000001",
47343 => "0000000000000001",47344 => "0000000000000001",
47345 => "0000000000000001",47346 => "0000000000000001",
47347 => "0000000000000001",47348 => "0000000000000001",
47349 => "0000000000000001",47350 => "0000000000000001",
47351 => "0000000000000001",47352 => "0000000000000001",
47353 => "0000000000000001",47354 => "0000000000000001",
47355 => "0000000000000001",47356 => "0000000000000001",
47357 => "0000000000000001",47358 => "0000000000000001",
47359 => "0000000000000001",47360 => "0000000000000001",
47361 => "0000000000000001",47362 => "0000000000000001",
47363 => "0000000000000001",47364 => "0000000000000001",
47365 => "0000000000000001",47366 => "0000000000000001",
47367 => "0000000000000001",47368 => "0000000000000001",
47369 => "0000000000000001",47370 => "0000000000000001",
47371 => "0000000000000001",47372 => "0000000000000001",
47373 => "0000000000000001",47374 => "0000000000000001",
47375 => "0000000000000001",47376 => "0000000000000001",
47377 => "0000000000000001",47378 => "0000000000000001",
47379 => "0000000000000001",47380 => "0000000000000001",
47381 => "0000000000000001",47382 => "0000000000000001",
47383 => "0000000000000001",47384 => "0000000000000001",
47385 => "0000000000000001",47386 => "0000000000000001",
47387 => "0000000000000001",47388 => "0000000000000001",
47389 => "0000000000000001",47390 => "0000000000000001",
47391 => "0000000000000001",47392 => "0000000000000001",
47393 => "0000000000000001",47394 => "0000000000000001",
47395 => "0000000000000001",47396 => "0000000000000001",
47397 => "0000000000000001",47398 => "0000000000000001",
47399 => "0000000000000001",47400 => "0000000000000001",
47401 => "0000000000000001",47402 => "0000000000000001",
47403 => "0000000000000001",47404 => "0000000000000001",
47405 => "0000000000000001",47406 => "0000000000000001",
47407 => "0000000000000001",47408 => "0000000000000001",
47409 => "0000000000000001",47410 => "0000000000000001",
47411 => "0000000000000001",47412 => "0000000000000001",
47413 => "0000000000000001",47414 => "0000000000000001",
47415 => "0000000000000001",47416 => "0000000000000001",
47417 => "0000000000000001",47418 => "0000000000000001",
47419 => "0000000000000001",47420 => "0000000000000001",
47421 => "0000000000000001",47422 => "0000000000000001",
47423 => "0000000000000001",47424 => "0000000000000001",
47425 => "0000000000000001",47426 => "0000000000000001",
47427 => "0000000000000001",47428 => "0000000000000001",
47429 => "0000000000000001",47430 => "0000000000000001",
47431 => "0000000000000001",47432 => "0000000000000001",
47433 => "0000000000000001",47434 => "0000000000000001",
47435 => "0000000000000001",47436 => "0000000000000001",
47437 => "0000000000000001",47438 => "0000000000000001",
47439 => "0000000000000001",47440 => "0000000000000001",
47441 => "0000000000000001",47442 => "0000000000000001",
47443 => "0000000000000001",47444 => "0000000000000001",
47445 => "0000000000000001",47446 => "0000000000000001",
47447 => "0000000000000001",47448 => "0000000000000001",
47449 => "0000000000000001",47450 => "0000000000000001",
47451 => "0000000000000001",47452 => "0000000000000001",
47453 => "0000000000000001",47454 => "0000000000000001",
47455 => "0000000000000001",47456 => "0000000000000001",
47457 => "0000000000000001",47458 => "0000000000000001",
47459 => "0000000000000001",47460 => "0000000000000001",
47461 => "0000000000000001",47462 => "0000000000000001",
47463 => "0000000000000001",47464 => "0000000000000001",
47465 => "0000000000000001",47466 => "0000000000000001",
47467 => "0000000000000001",47468 => "0000000000000001",
47469 => "0000000000000001",47470 => "0000000000000001",
47471 => "0000000000000001",47472 => "0000000000000001",
47473 => "0000000000000001",47474 => "0000000000000001",
47475 => "0000000000000001",47476 => "0000000000000001",
47477 => "0000000000000001",47478 => "0000000000000001",
47479 => "0000000000000001",47480 => "0000000000000001",
47481 => "0000000000000001",47482 => "0000000000000001",
47483 => "0000000000000001",47484 => "0000000000000001",
47485 => "0000000000000001",47486 => "0000000000000001",
47487 => "0000000000000001",47488 => "0000000000000001",
47489 => "0000000000000001",47490 => "0000000000000001",
47491 => "0000000000000001",47492 => "0000000000000001",
47493 => "0000000000000001",47494 => "0000000000000001",
47495 => "0000000000000001",47496 => "0000000000000001",
47497 => "0000000000000001",47498 => "0000000000000001",
47499 => "0000000000000001",47500 => "0000000000000001",
47501 => "0000000000000001",47502 => "0000000000000001",
47503 => "0000000000000001",47504 => "0000000000000001",
47505 => "0000000000000001",47506 => "0000000000000001",
47507 => "0000000000000001",47508 => "0000000000000001",
47509 => "0000000000000001",47510 => "0000000000000001",
47511 => "0000000000000001",47512 => "0000000000000001",
47513 => "0000000000000001",47514 => "0000000000000001",
47515 => "0000000000000001",47516 => "0000000000000001",
47517 => "0000000000000001",47518 => "0000000000000001",
47519 => "0000000000000001",47520 => "0000000000000001",
47521 => "0000000000000001",47522 => "0000000000000001",
47523 => "0000000000000001",47524 => "0000000000000001",
47525 => "0000000000000001",47526 => "0000000000000001",
47527 => "0000000000000001",47528 => "0000000000000001",
47529 => "0000000000000001",47530 => "0000000000000001",
47531 => "0000000000000001",47532 => "0000000000000001",
47533 => "0000000000000001",47534 => "0000000000000001",
47535 => "0000000000000001",47536 => "0000000000000001",
47537 => "0000000000000001",47538 => "0000000000000001",
47539 => "0000000000000001",47540 => "0000000000000001",
47541 => "0000000000000001",47542 => "0000000000000001",
47543 => "0000000000000001",47544 => "0000000000000001",
47545 => "0000000000000001",47546 => "0000000000000001",
47547 => "0000000000000001",47548 => "0000000000000001",
47549 => "0000000000000001",47550 => "0000000000000001",
47551 => "0000000000000001",47552 => "0000000000000001",
47553 => "0000000000000001",47554 => "0000000000000001",
47555 => "0000000000000001",47556 => "0000000000000001",
47557 => "0000000000000001",47558 => "0000000000000001",
47559 => "0000000000000001",47560 => "0000000000000001",
47561 => "0000000000000001",47562 => "0000000000000001",
47563 => "0000000000000001",47564 => "0000000000000001",
47565 => "0000000000000001",47566 => "0000000000000001",
47567 => "0000000000000001",47568 => "0000000000000001",
47569 => "0000000000000001",47570 => "0000000000000001",
47571 => "0000000000000001",47572 => "0000000000000001",
47573 => "0000000000000001",47574 => "0000000000000001",
47575 => "0000000000000001",47576 => "0000000000000001",
47577 => "0000000000000001",47578 => "0000000000000001",
47579 => "0000000000000001",47580 => "0000000000000001",
47581 => "0000000000000001",47582 => "0000000000000001",
47583 => "0000000000000001",47584 => "0000000000000001",
47585 => "0000000000000001",47586 => "0000000000000001",
47587 => "0000000000000001",47588 => "0000000000000001",
47589 => "0000000000000001",47590 => "0000000000000001",
47591 => "0000000000000001",47592 => "0000000000000001",
47593 => "0000000000000001",47594 => "0000000000000001",
47595 => "0000000000000001",47596 => "0000000000000001",
47597 => "0000000000000001",47598 => "0000000000000001",
47599 => "0000000000000001",47600 => "0000000000000001",
47601 => "0000000000000001",47602 => "0000000000000001",
47603 => "0000000000000001",47604 => "0000000000000001",
47605 => "0000000000000001",47606 => "0000000000000001",
47607 => "0000000000000001",47608 => "0000000000000001",
47609 => "0000000000000001",47610 => "0000000000000001",
47611 => "0000000000000001",47612 => "0000000000000001",
47613 => "0000000000000001",47614 => "0000000000000001",
47615 => "0000000000000001",47616 => "0000000000000001",
47617 => "0000000000000001",47618 => "0000000000000001",
47619 => "0000000000000001",47620 => "0000000000000001",
47621 => "0000000000000001",47622 => "0000000000000001",
47623 => "0000000000000001",47624 => "0000000000000001",
47625 => "0000000000000001",47626 => "0000000000000001",
47627 => "0000000000000001",47628 => "0000000000000001",
47629 => "0000000000000001",47630 => "0000000000000001",
47631 => "0000000000000001",47632 => "0000000000000001",
47633 => "0000000000000001",47634 => "0000000000000001",
47635 => "0000000000000001",47636 => "0000000000000001",
47637 => "0000000000000001",47638 => "0000000000000001",
47639 => "0000000000000001",47640 => "0000000000000001",
47641 => "0000000000000001",47642 => "0000000000000001",
47643 => "0000000000000001",47644 => "0000000000000001",
47645 => "0000000000000001",47646 => "0000000000000001",
47647 => "0000000000000001",47648 => "0000000000000001",
47649 => "0000000000000001",47650 => "0000000000000001",
47651 => "0000000000000001",47652 => "0000000000000001",
47653 => "0000000000000001",47654 => "0000000000000001",
47655 => "0000000000000001",47656 => "0000000000000001",
47657 => "0000000000000001",47658 => "0000000000000001",
47659 => "0000000000000001",47660 => "0000000000000001",
47661 => "0000000000000001",47662 => "0000000000000001",
47663 => "0000000000000001",47664 => "0000000000000001",
47665 => "0000000000000001",47666 => "0000000000000001",
47667 => "0000000000000001",47668 => "0000000000000001",
47669 => "0000000000000001",47670 => "0000000000000001",
47671 => "0000000000000001",47672 => "0000000000000001",
47673 => "0000000000000001",47674 => "0000000000000001",
47675 => "0000000000000001",47676 => "0000000000000001",
47677 => "0000000000000001",47678 => "0000000000000001",
47679 => "0000000000000001",47680 => "0000000000000001",
47681 => "0000000000000001",47682 => "0000000000000001",
47683 => "0000000000000001",47684 => "0000000000000001",
47685 => "0000000000000001",47686 => "0000000000000001",
47687 => "0000000000000001",47688 => "0000000000000001",
47689 => "0000000000000001",47690 => "0000000000000001",
47691 => "0000000000000001",47692 => "0000000000000001",
47693 => "0000000000000001",47694 => "0000000000000001",
47695 => "0000000000000001",47696 => "0000000000000001",
47697 => "0000000000000001",47698 => "0000000000000001",
47699 => "0000000000000001",47700 => "0000000000000001",
47701 => "0000000000000001",47702 => "0000000000000001",
47703 => "0000000000000001",47704 => "0000000000000001",
47705 => "0000000000000000",47706 => "0000000000000000",
47707 => "0000000000000000",47708 => "0000000000000000",
47709 => "0000000000000000",47710 => "0000000000000000",
47711 => "0000000000000000",47712 => "0000000000000000",
47713 => "0000000000000000",47714 => "0000000000000000",
47715 => "0000000000000000",47716 => "0000000000000000",
47717 => "0000000000000000",47718 => "0000000000000000",
47719 => "0000000000000000",47720 => "0000000000000000",
47721 => "0000000000000000",47722 => "0000000000000000",
47723 => "0000000000000000",47724 => "0000000000000000",
47725 => "0000000000000000",47726 => "0000000000000000",
47727 => "0000000000000000",47728 => "0000000000000000",
47729 => "0000000000000000",47730 => "0000000000000000",
47731 => "0000000000000000",47732 => "0000000000000000",
47733 => "0000000000000000",47734 => "0000000000000000",
47735 => "0000000000000000",47736 => "0000000000000000",
47737 => "0000000000000000",47738 => "0000000000000000",
47739 => "0000000000000000",47740 => "0000000000000000",
47741 => "0000000000000000",47742 => "0000000000000000",
47743 => "0000000000000000",47744 => "0000000000000000",
47745 => "0000000000000000",47746 => "0000000000000000",
47747 => "0000000000000000",47748 => "0000000000000000",
47749 => "0000000000000000",47750 => "0000000000000000",
47751 => "0000000000000000",47752 => "0000000000000000",
47753 => "0000000000000000",47754 => "0000000000000000",
47755 => "0000000000000000",47756 => "0000000000000000",
47757 => "0000000000000000",47758 => "0000000000000000",
47759 => "0000000000000000",47760 => "0000000000000000",
47761 => "0000000000000000",47762 => "0000000000000000",
47763 => "0000000000000000",47764 => "0000000000000000",
47765 => "0000000000000000",47766 => "0000000000000000",
47767 => "0000000000000000",47768 => "0000000000000000",
47769 => "0000000000000000",47770 => "0000000000000000",
47771 => "0000000000000000",47772 => "0000000000000000",
47773 => "0000000000000000",47774 => "0000000000000000",
47775 => "0000000000000000",47776 => "0000000000000000",
47777 => "0000000000000000",47778 => "0000000000000000",
47779 => "0000000000000000",47780 => "0000000000000000",
47781 => "0000000000000000",47782 => "0000000000000000",
47783 => "0000000000000000",47784 => "0000000000000000",
47785 => "0000000000000000",47786 => "0000000000000000",
47787 => "0000000000000000",47788 => "0000000000000000",
47789 => "0000000000000000",47790 => "0000000000000000",
47791 => "0000000000000000",47792 => "0000000000000000",
47793 => "0000000000000000",47794 => "0000000000000000",
47795 => "0000000000000000",47796 => "0000000000000000",
47797 => "0000000000000000",47798 => "0000000000000000",
47799 => "0000000000000000",47800 => "0000000000000000",
47801 => "0000000000000000",47802 => "0000000000000000",
47803 => "0000000000000000",47804 => "0000000000000000",
47805 => "0000000000000000",47806 => "0000000000000000",
47807 => "0000000000000000",47808 => "0000000000000000",
47809 => "0000000000000000",47810 => "0000000000000000",
47811 => "0000000000000000",47812 => "0000000000000000",
47813 => "0000000000000000",47814 => "0000000000000000",
47815 => "0000000000000000",47816 => "0000000000000000",
47817 => "0000000000000000",47818 => "0000000000000000",
47819 => "0000000000000000",47820 => "0000000000000000",
47821 => "0000000000000000",47822 => "0000000000000000",
47823 => "0000000000000000",47824 => "0000000000000000",
47825 => "0000000000000000",47826 => "0000000000000000",
47827 => "0000000000000000",47828 => "0000000000000000",
47829 => "0000000000000000",47830 => "0000000000000000",
47831 => "0000000000000000",47832 => "0000000000000000",
47833 => "0000000000000000",47834 => "0000000000000000",
47835 => "0000000000000000",47836 => "0000000000000000",
47837 => "0000000000000000",47838 => "0000000000000000",
47839 => "0000000000000000",47840 => "0000000000000000",
47841 => "0000000000000000",47842 => "0000000000000000",
47843 => "0000000000000000",47844 => "0000000000000000",
47845 => "0000000000000000",47846 => "0000000000000000",
47847 => "0000000000000000",47848 => "0000000000000000",
47849 => "0000000000000000",47850 => "0000000000000000",
47851 => "0000000000000000",47852 => "0000000000000000",
47853 => "0000000000000000",47854 => "0000000000000000",
47855 => "0000000000000000",47856 => "0000000000000000",
47857 => "0000000000000000",47858 => "0000000000000000",
47859 => "0000000000000000",47860 => "0000000000000000",
47861 => "0000000000000000",47862 => "0000000000000000",
47863 => "0000000000000000",47864 => "0000000000000000",
47865 => "0000000000000000",47866 => "0000000000000000",
47867 => "0000000000000000",47868 => "0000000000000000",
47869 => "0000000000000000",47870 => "0000000000000000",
47871 => "0000000000000000",47872 => "0000000000000000",
47873 => "0000000000000000",47874 => "0000000000000000",
47875 => "0000000000000000",47876 => "0000000000000000",
47877 => "0000000000000000",47878 => "0000000000000000",
47879 => "0000000000000000",47880 => "0000000000000000",
47881 => "0000000000000000",47882 => "0000000000000000",
47883 => "0000000000000000",47884 => "0000000000000000",
47885 => "0000000000000000",47886 => "0000000000000000",
47887 => "0000000000000000",47888 => "0000000000000000",
47889 => "0000000000000000",47890 => "0000000000000000",
47891 => "0000000000000000",47892 => "0000000000000000",
47893 => "0000000000000000",47894 => "0000000000000000",
47895 => "0000000000000000",47896 => "0000000000000000",
47897 => "0000000000000000",47898 => "0000000000000000",
47899 => "0000000000000000",47900 => "0000000000000000",
47901 => "0000000000000000",47902 => "0000000000000000",
47903 => "0000000000000000",47904 => "0000000000000000",
47905 => "0000000000000000",47906 => "0000000000000000",
47907 => "0000000000000000",47908 => "0000000000000000",
47909 => "0000000000000000",47910 => "0000000000000000",
47911 => "0000000000000000",47912 => "0000000000000000",
47913 => "0000000000000000",47914 => "0000000000000000",
47915 => "0000000000000000",47916 => "0000000000000000",
47917 => "0000000000000000",47918 => "0000000000000000",
47919 => "0000000000000000",47920 => "0000000000000000",
47921 => "0000000000000000",47922 => "0000000000000000",
47923 => "0000000000000000",47924 => "0000000000000000",
47925 => "0000000000000000",47926 => "0000000000000000",
47927 => "0000000000000000",47928 => "0000000000000000",
47929 => "0000000000000000",47930 => "0000000000000000",
47931 => "0000000000000000",47932 => "0000000000000000",
47933 => "0000000000000000",47934 => "0000000000000000",
47935 => "0000000000000000",47936 => "0000000000000000",
47937 => "0000000000000000",47938 => "0000000000000000",
47939 => "0000000000000000",47940 => "0000000000000000",
47941 => "0000000000000000",47942 => "0000000000000000",
47943 => "0000000000000000",47944 => "0000000000000000",
47945 => "0000000000000000",47946 => "0000000000000000",
47947 => "0000000000000000",47948 => "0000000000000000",
47949 => "0000000000000000",47950 => "0000000000000000",
47951 => "0000000000000000",47952 => "0000000000000000",
47953 => "0000000000000000",47954 => "0000000000000000",
47955 => "0000000000000000",47956 => "0000000000000000",
47957 => "0000000000000000",47958 => "0000000000000000",
47959 => "0000000000000000",47960 => "0000000000000000",
47961 => "0000000000000000",47962 => "0000000000000000",
47963 => "0000000000000000",47964 => "0000000000000000",
47965 => "0000000000000000",47966 => "0000000000000000",
47967 => "0000000000000000",47968 => "0000000000000000",
47969 => "0000000000000000",47970 => "0000000000000000",
47971 => "0000000000000000",47972 => "0000000000000000",
47973 => "0000000000000000",47974 => "0000000000000000",
47975 => "0000000000000000",47976 => "0000000000000000",
47977 => "0000000000000000",47978 => "0000000000000000",
47979 => "0000000000000000",47980 => "0000000000000000",
47981 => "0000000000000000",47982 => "0000000000000000",
47983 => "0000000000000000",47984 => "0000000000000000",
47985 => "0000000000000000",47986 => "0000000000000000",
47987 => "0000000000000000",47988 => "0000000000000000",
47989 => "0000000000000000",47990 => "0000000000000000",
47991 => "0000000000000000",47992 => "0000000000000000",
47993 => "0000000000000000",47994 => "0000000000000000",
47995 => "0000000000000000",47996 => "0000000000000000",
47997 => "0000000000000000",47998 => "0000000000000000",
47999 => "0000000000000000",48000 => "0000000000000000",
48001 => "0000000000000000",48002 => "0000000000000000",
48003 => "0000000000000000",48004 => "0000000000000000",
48005 => "0000000000000000",48006 => "0000000000000000",
48007 => "0000000000000000",48008 => "0000000000000000",
48009 => "0000000000000000",48010 => "0000000000000000",
48011 => "0000000000000000",48012 => "0000000000000000",
48013 => "0000000000000000",48014 => "0000000000000000",
48015 => "0000000000000000",48016 => "0000000000000000",
48017 => "0000000000000000",48018 => "0000000000000000",
48019 => "0000000000000000",48020 => "0000000000000000",
48021 => "0000000000000000",48022 => "0000000000000000",
48023 => "0000000000000000",48024 => "0000000000000000",
48025 => "0000000000000000",48026 => "0000000000000000",
48027 => "0000000000000000",48028 => "0000000000000000",
48029 => "0000000000000000",48030 => "0000000000000000",
48031 => "0000000000000000",48032 => "0000000000000000",
48033 => "0000000000000000",48034 => "0000000000000000",
48035 => "0000000000000000",48036 => "0000000000000000",
48037 => "0000000000000000",48038 => "0000000000000000",
48039 => "0000000000000000",48040 => "0000000000000000",
48041 => "0000000000000000",48042 => "0000000000000000",
48043 => "0000000000000000",48044 => "0000000000000000",
48045 => "0000000000000000",48046 => "0000000000000000",
48047 => "0000000000000000",48048 => "0000000000000000",
48049 => "0000000000000000",48050 => "0000000000000000",
48051 => "0000000000000000",48052 => "0000000000000000",
48053 => "0000000000000000",48054 => "0000000000000000",
48055 => "0000000000000000",48056 => "0000000000000000",
48057 => "0000000000000000",48058 => "0000000000000000",
48059 => "0000000000000000",48060 => "0000000000000000",
48061 => "0000000000000000",48062 => "0000000000000000",
48063 => "0000000000000000",48064 => "0000000000000000",
48065 => "0000000000000000",48066 => "0000000000000000",
48067 => "0000000000000000",48068 => "0000000000000000",
48069 => "0000000000000000",48070 => "0000000000000000",
48071 => "0000000000000000",48072 => "0000000000000000",
48073 => "0000000000000000",48074 => "0000000000000000",
48075 => "0000000000000000",48076 => "0000000000000000",
48077 => "0000000000000000",48078 => "0000000000000000",
48079 => "0000000000000000",48080 => "0000000000000000",
48081 => "0000000000000000",48082 => "0000000000000000",
48083 => "0000000000000000",48084 => "0000000000000000",
48085 => "0000000000000000",48086 => "0000000000000000",
48087 => "0000000000000000",48088 => "0000000000000000",
48089 => "0000000000000000",48090 => "0000000000000000",
48091 => "0000000000000000",48092 => "0000000000000000",
48093 => "0000000000000000",48094 => "0000000000000000",
48095 => "0000000000000000",48096 => "0000000000000000",
48097 => "0000000000000000",48098 => "0000000000000000",
48099 => "0000000000000000",48100 => "0000000000000000",
48101 => "0000000000000000",48102 => "0000000000000000",
48103 => "0000000000000000",48104 => "0000000000000001",
48105 => "0000000000000001",48106 => "0000000000000001",
48107 => "0000000000000001",48108 => "0000000000000001",
48109 => "0000000000000001",48110 => "0000000000000001",
48111 => "0000000000000001",48112 => "0000000000000001",
48113 => "0000000000000001",48114 => "0000000000000001",
48115 => "0000000000000001",48116 => "0000000000000001",
48117 => "0000000000000001",48118 => "0000000000000001",
48119 => "0000000000000001",48120 => "0000000000000001",
48121 => "0000000000000001",48122 => "0000000000000001",
48123 => "0000000000000001",48124 => "0000000000000001",
48125 => "0000000000000001",48126 => "0000000000000001",
48127 => "0000000000000001",48128 => "0000000000000001",
48129 => "0000000000000001",48130 => "0000000000000001",
48131 => "0000000000000001",48132 => "0000000000000001",
48133 => "0000000000000001",48134 => "0000000000000001",
48135 => "0000000000000001",48136 => "0000000000000001",
48137 => "0000000000000001",48138 => "0000000000000001",
48139 => "0000000000000001",48140 => "0000000000000001",
48141 => "0000000000000001",48142 => "0000000000000001",
48143 => "0000000000000001",48144 => "0000000000000001",
48145 => "0000000000000001",48146 => "0000000000000001",
48147 => "0000000000000001",48148 => "0000000000000001",
48149 => "0000000000000001",48150 => "0000000000000001",
48151 => "0000000000000001",48152 => "0000000000000001",
48153 => "0000000000000001",48154 => "0000000000000001",
48155 => "0000000000000001",48156 => "0000000000000001",
48157 => "0000000000000001",48158 => "0000000000000001",
48159 => "0000000000000001",48160 => "0000000000000001",
48161 => "0000000000000001",48162 => "0000000000000001",
48163 => "0000000000000001",48164 => "0000000000000001",
48165 => "0000000000000001",48166 => "0000000000000001",
48167 => "0000000000000001",48168 => "0000000000000001",
48169 => "0000000000000001",48170 => "0000000000000001",
48171 => "0000000000000001",48172 => "0000000000000001",
48173 => "0000000000000001",48174 => "0000000000000001",
48175 => "0000000000000001",48176 => "0000000000000001",
48177 => "0000000000000001",48178 => "0000000000000001",
48179 => "0000000000000001",48180 => "0000000000000001",
48181 => "0000000000000001",48182 => "0000000000000001",
48183 => "0000000000000001",48184 => "0000000000000001",
48185 => "0000000000000001",48186 => "0000000000000001",
48187 => "0000000000000001",48188 => "0000000000000001",
48189 => "0000000000000001",48190 => "0000000000000001",
48191 => "0000000000000001",48192 => "0000000000000001",
48193 => "0000000000000001",48194 => "0000000000000001",
48195 => "0000000000000001",48196 => "0000000000000001",
48197 => "0000000000000001",48198 => "0000000000000001",
48199 => "0000000000000001",48200 => "0000000000000001",
48201 => "0000000000000001",48202 => "0000000000000001",
48203 => "0000000000000001",48204 => "0000000000000001",
48205 => "0000000000000001",48206 => "0000000000000001",
48207 => "0000000000000001",48208 => "0000000000000001",
48209 => "0000000000000001",48210 => "0000000000000001",
48211 => "0000000000000001",48212 => "0000000000000001",
48213 => "0000000000000001",48214 => "0000000000000001",
48215 => "0000000000000001",48216 => "0000000000000001",
48217 => "0000000000000001",48218 => "0000000000000001",
48219 => "0000000000000001",48220 => "0000000000000001",
48221 => "0000000000000001",48222 => "0000000000000001",
48223 => "0000000000000001",48224 => "0000000000000001",
48225 => "0000000000000001",48226 => "0000000000000001",
48227 => "0000000000000001",48228 => "0000000000000001",
48229 => "0000000000000001",48230 => "0000000000000001",
48231 => "0000000000000001",48232 => "0000000000000001",
48233 => "0000000000000001",48234 => "0000000000000001",
48235 => "0000000000000001",48236 => "0000000000000001",
48237 => "0000000000000001",48238 => "0000000000000001",
48239 => "0000000000000001",48240 => "0000000000000001",
48241 => "0000000000000001",48242 => "0000000000000001",
48243 => "0000000000000001",48244 => "0000000000000001",
48245 => "0000000000000001",48246 => "0000000000000001",
48247 => "0000000000000001",48248 => "0000000000000001",
48249 => "0000000000000001",48250 => "0000000000000001",
48251 => "0000000000000001",48252 => "0000000000000001",
48253 => "0000000000000001",48254 => "0000000000000001",
48255 => "0000000000000001",48256 => "0000000000000001",
48257 => "0000000000000001",48258 => "0000000000000001",
48259 => "0000000000000001",48260 => "0000000000000001",
48261 => "0000000000000001",48262 => "0000000000000001",
48263 => "0000000000000001",48264 => "0000000000000001",
48265 => "0000000000000001",48266 => "0000000000000001",
48267 => "0000000000000001",48268 => "0000000000000001",
48269 => "0000000000000001",48270 => "0000000000000001",
48271 => "0000000000000001",48272 => "0000000000000001",
48273 => "0000000000000001",48274 => "0000000000000001",
48275 => "0000000000000001",48276 => "0000000000000001",
48277 => "0000000000000001",48278 => "0000000000000001",
48279 => "0000000000000001",48280 => "0000000000000001",
48281 => "0000000000000001",48282 => "0000000000000001",
48283 => "0000000000000001",48284 => "0000000000000001",
48285 => "0000000000000001",48286 => "0000000000000001",
48287 => "0000000000000001",48288 => "0000000000000001",
48289 => "0000000000000001",48290 => "0000000000000001",
48291 => "0000000000000001",48292 => "0000000000000001",
48293 => "0000000000000001",48294 => "0000000000000001",
48295 => "0000000000000001",48296 => "0000000000000001",
48297 => "0000000000000001",48298 => "0000000000000001",
48299 => "0000000000000001",48300 => "0000000000000001",
48301 => "0000000000000001",48302 => "0000000000000001",
48303 => "0000000000000001",48304 => "0000000000000001",
48305 => "0000000000000001",48306 => "0000000000000001",
48307 => "0000000000000001",48308 => "0000000000000001",
48309 => "0000000000000001",48310 => "0000000000000001",
48311 => "0000000000000001",48312 => "0000000000000001",
48313 => "0000000000000001",48314 => "0000000000000001",
48315 => "0000000000000001",48316 => "0000000000000001",
48317 => "0000000000000001",48318 => "0000000000000001",
48319 => "0000000000000001",48320 => "0000000000000001",
48321 => "0000000000000001",48322 => "0000000000000001",
48323 => "0000000000000001",48324 => "0000000000000001",
48325 => "0000000000000001",48326 => "0000000000000001",
48327 => "0000000000000001",48328 => "0000000000000001",
48329 => "0000000000000001",48330 => "0000000000000001",
48331 => "0000000000000001",48332 => "0000000000000001",
48333 => "0000000000000001",48334 => "0000000000000001",
48335 => "0000000000000001",48336 => "0000000000000001",
48337 => "0000000000000001",48338 => "0000000000000001",
48339 => "0000000000000001",48340 => "0000000000000001",
48341 => "0000000000000001",48342 => "0000000000000001",
48343 => "0000000000000001",48344 => "0000000000000001",
48345 => "0000000000000001",48346 => "0000000000000001",
48347 => "0000000000000001",48348 => "0000000000000001",
48349 => "0000000000000001",48350 => "0000000000000001",
48351 => "0000000000000001",48352 => "0000000000000001",
48353 => "0000000000000001",48354 => "0000000000000001",
48355 => "0000000000000001",48356 => "0000000000000001",
48357 => "0000000000000001",48358 => "0000000000000001",
48359 => "0000000000000001",48360 => "0000000000000001",
48361 => "0000000000000001",48362 => "0000000000000001",
48363 => "0000000000000001",48364 => "0000000000000001",
48365 => "0000000000000001",48366 => "0000000000000001",
48367 => "0000000000000001",48368 => "0000000000000001",
48369 => "0000000000000001",48370 => "0000000000000001",
48371 => "0000000000000001",48372 => "0000000000000001",
48373 => "0000000000000001",48374 => "0000000000000001",
48375 => "0000000000000001",48376 => "0000000000000001",
48377 => "0000000000000001",48378 => "0000000000000001",
48379 => "0000000000000001",48380 => "0000000000000001",
48381 => "0000000000000001",48382 => "0000000000000001",
48383 => "0000000000000001",48384 => "0000000000000001",
48385 => "0000000000000001",48386 => "0000000000000001",
48387 => "0000000000000001",48388 => "0000000000000001",
48389 => "0000000000000001",48390 => "0000000000000001",
48391 => "0000000000000001",48392 => "0000000000000001",
48393 => "0000000000000001",48394 => "0000000000000001",
48395 => "0000000000000001",48396 => "0000000000000001",
48397 => "0000000000000001",48398 => "0000000000000001",
48399 => "0000000000000001",48400 => "0000000000000001",
48401 => "0000000000000001",48402 => "0000000000000001",
48403 => "0000000000000001",48404 => "0000000000000001",
48405 => "0000000000000001",48406 => "0000000000000001",
48407 => "0000000000000001",48408 => "0000000000000001",
48409 => "0000000000000001",48410 => "0000000000000001",
48411 => "0000000000000001",48412 => "0000000000000001",
48413 => "0000000000000001",48414 => "0000000000000001",
48415 => "0000000000000001",48416 => "0000000000000001",
48417 => "0000000000000001",48418 => "0000000000000001",
48419 => "0000000000000001",48420 => "0000000000000001",
48421 => "0000000000000001",48422 => "0000000000000001",
48423 => "0000000000000001",48424 => "0000000000000001",
48425 => "0000000000000001",48426 => "0000000000000001",
48427 => "0000000000000001",48428 => "0000000000000001",
48429 => "0000000000000001",48430 => "0000000000000001",
48431 => "0000000000000001",48432 => "0000000000000001",
48433 => "0000000000000001",48434 => "0000000000000001",
48435 => "0000000000000001",48436 => "0000000000000001",
48437 => "0000000000000001",48438 => "0000000000000001",
48439 => "0000000000000001",48440 => "0000000000000001",
48441 => "0000000000000001",48442 => "0000000000000001",
48443 => "0000000000000001",48444 => "0000000000000001",
48445 => "0000000000000001",48446 => "0000000000000001",
48447 => "0000000000000001",48448 => "0000000000000001",
48449 => "0000000000000001",48450 => "0000000000000001",
48451 => "0000000000000001",48452 => "0000000000000001",
48453 => "0000000000000001",48454 => "0000000000000001",
48455 => "0000000000000001",48456 => "0000000000000001",
48457 => "0000000000000001",48458 => "0000000000000001",
48459 => "0000000000000001",48460 => "0000000000000001",
48461 => "0000000000000001",48462 => "0000000000000001",
48463 => "0000000000000001",48464 => "0000000000000001",
48465 => "0000000000000001",48466 => "0000000000000001",
48467 => "0000000000000001",48468 => "0000000000000001",
48469 => "0000000000000001",48470 => "0000000000000001",
48471 => "0000000000000001",48472 => "0000000000000001",
48473 => "0000000000000001",48474 => "0000000000000001",
48475 => "0000000000000001",48476 => "0000000000000001",
48477 => "0000000000000001",48478 => "0000000000000001",
48479 => "0000000000000001",48480 => "0000000000000001",
48481 => "0000000000000001",48482 => "0000000000000001",
48483 => "0000000000000001",48484 => "0000000000000001",
48485 => "0000000000000001",48486 => "0000000000000001",
48487 => "0000000000000001",48488 => "0000000000000001",
48489 => "0000000000000001",48490 => "0000000000000001",
48491 => "0000000000000001",48492 => "0000000000000001",
48493 => "0000000000000001",48494 => "0000000000000001",
48495 => "0000000000000001",48496 => "0000000000000001",
48497 => "0000000000000001",48498 => "0000000000000001",
48499 => "0000000000000001",48500 => "0000000000000001",
48501 => "0000000000000001",48502 => "0000000000000001",
48503 => "0000000000000001",48504 => "0000000000000001",
48505 => "0000000000000001",48506 => "0000000000000001",
48507 => "0000000000000001",48508 => "0000000000000001",
48509 => "0000000000000001",48510 => "0000000000000001",
48511 => "0000000000000001",48512 => "0000000000000001",
48513 => "0000000000000001",48514 => "0000000000000001",
48515 => "0000000000000001",48516 => "0000000000000001",
48517 => "0000000000000001",48518 => "0000000000000001",
48519 => "0000000000000001",48520 => "0000000000000001",
48521 => "0000000000000001",48522 => "0000000000000001",
48523 => "0000000000000001",48524 => "0000000000000001",
48525 => "0000000000000001",48526 => "0000000000000001",
48527 => "0000000000000001",48528 => "0000000000000001",
48529 => "0000000000000001",48530 => "0000000000000001",
48531 => "0000000000000001",48532 => "0000000000000001",
48533 => "0000000000000001",48534 => "0000000000000001",
48535 => "0000000000000001",48536 => "0000000000000001",
48537 => "0000000000000001",48538 => "0000000000000001",
48539 => "0000000000000001",48540 => "0000000000000001",
48541 => "0000000000000001",48542 => "0000000000000001",
48543 => "0000000000000001",48544 => "0000000000000001",
48545 => "0000000000000001",48546 => "0000000000000001",
48547 => "0000000000000001",48548 => "0000000000000001",
48549 => "0000000000000001",48550 => "0000000000000001",
48551 => "0000000000000001",48552 => "0000000000000001",
48553 => "0000000000000001",48554 => "0000000000000001",
48555 => "0000000000000001",48556 => "0000000000000001",
48557 => "0000000000000001",48558 => "0000000000000001",
48559 => "0000000000000001",48560 => "0000000000000001",
48561 => "0000000000000001",48562 => "0000000000000001",
48563 => "0000000000000001",48564 => "0000000000000001",
48565 => "0000000000000001",48566 => "0000000000000001",
48567 => "0000000000000001",48568 => "0000000000000001",
48569 => "0000000000000001",48570 => "0000000000000001",
48571 => "0000000000000001",48572 => "0000000000000001",
48573 => "0000000000000001",48574 => "0000000000000001",
48575 => "0000000000000001",48576 => "0000000000000001",
48577 => "0000000000000001",48578 => "0000000000000001",
48579 => "0000000000000001",48580 => "0000000000000001",
48581 => "0000000000000001",48582 => "0000000000000001",
48583 => "0000000000000001",48584 => "0000000000000001",
48585 => "0000000000000001",48586 => "0000000000000001",
48587 => "0000000000000001",48588 => "0000000000000001",
48589 => "0000000000000001",48590 => "0000000000000001",
48591 => "0000000000000001",48592 => "0000000000000001",
48593 => "0000000000000001",48594 => "0000000000000001",
48595 => "0000000000000001",48596 => "0000000000000001",
48597 => "0000000000000001",48598 => "0000000000000001",
48599 => "0000000000000001",48600 => "0000000000000001",
48601 => "0000000000000001",48602 => "0000000000000001",
48603 => "0000000000000001",48604 => "0000000000000001",
48605 => "0000000000000001",48606 => "0000000000000001",
48607 => "0000000000000001",48608 => "0000000000000001",
48609 => "0000000000000001",48610 => "0000000000000001",
48611 => "0000000000000001",48612 => "0000000000000001",
48613 => "0000000000000001",48614 => "0000000000000001",
48615 => "0000000000000001",48616 => "0000000000000001",
48617 => "0000000000000001",48618 => "0000000000000001",
48619 => "0000000000000001",48620 => "0000000000000001",
48621 => "0000000000000001",48622 => "0000000000000001",
48623 => "0000000000000001",48624 => "0000000000000001",
48625 => "0000000000000001",48626 => "0000000000000001",
48627 => "0000000000000001",48628 => "0000000000000001",
48629 => "0000000000000001",48630 => "0000000000000001",
48631 => "0000000000000001",48632 => "0000000000000001",
48633 => "0000000000000001",48634 => "0000000000000001",
48635 => "0000000000000001",48636 => "0000000000000001",
48637 => "0000000000000001",48638 => "0000000000000001",
48639 => "0000000000000001",48640 => "0000000000000001",
48641 => "0000000000000001",48642 => "0000000000000001",
48643 => "0000000000000001",48644 => "0000000000000001",
48645 => "0000000000000001",48646 => "0000000000000001",
48647 => "0000000000000001",48648 => "0000000000000001",
48649 => "0000000000000001",48650 => "0000000000000001",
48651 => "0000000000000001",48652 => "0000000000000001",
48653 => "0000000000000001",48654 => "0000000000000001",
48655 => "0000000000000001",48656 => "0000000000000001",
48657 => "0000000000000001",48658 => "0000000000000001",
48659 => "0000000000000001",48660 => "0000000000000001",
48661 => "0000000000000001",48662 => "0000000000000001",
48663 => "0000000000000001",48664 => "0000000000000001",
48665 => "0000000000000001",48666 => "0000000000000001",
48667 => "0000000000000001",48668 => "0000000000000001",
48669 => "0000000000000001",48670 => "0000000000000001",
48671 => "0000000000000001",48672 => "0000000000000001",
48673 => "0000000000000001",48674 => "0000000000000001",
48675 => "0000000000000001",48676 => "0000000000000001",
48677 => "0000000000000001",48678 => "0000000000000001",
48679 => "0000000000000001",48680 => "0000000000000001",
48681 => "0000000000000001",48682 => "0000000000000001",
48683 => "0000000000000001",48684 => "0000000000000001",
48685 => "0000000000000001",48686 => "0000000000000001",
48687 => "0000000000000001",48688 => "0000000000000001",
48689 => "0000000000000001",48690 => "0000000000000001",
48691 => "0000000000000001",48692 => "0000000000000001",
48693 => "0000000000000001",48694 => "0000000000000001",
48695 => "0000000000000001",48696 => "0000000000000001",
48697 => "0000000000000001",48698 => "0000000000000001",
48699 => "0000000000000001",48700 => "0000000000000001",
48701 => "0000000000000001",48702 => "0000000000000001",
48703 => "0000000000000001",48704 => "0000000000000001",
48705 => "0000000000000001",48706 => "0000000000000001",
48707 => "0000000000000001",48708 => "0000000000000001",
48709 => "0000000000000001",48710 => "0000000000000001",
48711 => "0000000000000001",48712 => "0000000000000001",
48713 => "0000000000000001",48714 => "0000000000000001",
48715 => "0000000000000001",48716 => "0000000000000001",
48717 => "0000000000000001",48718 => "0000000000000001",
48719 => "0000000000000001",48720 => "0000000000000001",
48721 => "0000000000000001",48722 => "0000000000000001",
48723 => "0000000000000001",48724 => "0000000000000001",
48725 => "0000000000000001",48726 => "0000000000000001",
48727 => "0000000000000001",48728 => "0000000000000001",
48729 => "0000000000000001",48730 => "0000000000000001",
48731 => "0000000000000001",48732 => "0000000000000001",
48733 => "0000000000000001",48734 => "0000000000000001",
48735 => "0000000000000001",48736 => "0000000000000001",
48737 => "0000000000000001",48738 => "0000000000000001",
48739 => "0000000000000001",48740 => "0000000000000001",
48741 => "0000000000000001",48742 => "0000000000000001",
48743 => "0000000000000001",48744 => "0000000000000001",
48745 => "0000000000000001",48746 => "0000000000000001",
48747 => "0000000000000001",48748 => "0000000000000001",
48749 => "0000000000000001",48750 => "0000000000000001",
48751 => "0000000000000001",48752 => "0000000000000001",
48753 => "0000000000000001",48754 => "0000000000000001",
48755 => "0000000000000001",48756 => "0000000000000001",
48757 => "0000000000000001",48758 => "0000000000000001",
48759 => "0000000000000001",48760 => "0000000000000001",
48761 => "0000000000000001",48762 => "0000000000000001",
48763 => "0000000000000001",48764 => "0000000000000001",
48765 => "0000000000000001",48766 => "0000000000000001",
48767 => "0000000000000001",48768 => "0000000000000001",
48769 => "0000000000000001",48770 => "0000000000000001",
48771 => "0000000000000001",48772 => "0000000000000001",
48773 => "0000000000000001",48774 => "0000000000000001",
48775 => "0000000000000001",48776 => "0000000000000001",
48777 => "0000000000000001",48778 => "0000000000000001",
48779 => "0000000000000001",48780 => "0000000000000001",
48781 => "0000000000000001",48782 => "0000000000000001",
48783 => "0000000000000001",48784 => "0000000000000001",
48785 => "0000000000000001",48786 => "0000000000000001",
48787 => "0000000000000001",48788 => "0000000000000001",
48789 => "0000000000000001",48790 => "0000000000000001",
48791 => "0000000000000001",48792 => "0000000000000001",
48793 => "0000000000000001",48794 => "0000000000000001",
48795 => "0000000000000001",48796 => "0000000000000001",
48797 => "0000000000000001",48798 => "0000000000000001",
48799 => "0000000000000001",48800 => "0000000000000001",
48801 => "0000000000000001",48802 => "0000000000000001",
48803 => "0000000000000001",48804 => "0000000000000001",
48805 => "0000000000000001",48806 => "0000000000000001",
48807 => "0000000000000001",48808 => "0000000000000001",
48809 => "0000000000000001",48810 => "0000000000000001",
48811 => "0000000000000001",48812 => "0000000000000001",
48813 => "0000000000000001",48814 => "0000000000000001",
48815 => "0000000000000001",48816 => "0000000000000001",
48817 => "0000000000000001",48818 => "0000000000000001",
48819 => "0000000000000001",48820 => "0000000000000001",
48821 => "0000000000000001",48822 => "0000000000000001",
48823 => "0000000000000001",48824 => "0000000000000001",
48825 => "0000000000000001",48826 => "0000000000000001",
48827 => "0000000000000001",48828 => "0000000000000001",
48829 => "0000000000000001",48830 => "0000000000000001",
48831 => "0000000000000001",48832 => "0000000000000001",
48833 => "0000000000000001",48834 => "0000000000000001",
48835 => "0000000000000001",48836 => "0000000000000001",
48837 => "0000000000000001",48838 => "0000000000000001",
48839 => "0000000000000001",48840 => "0000000000000001",
48841 => "0000000000000001",48842 => "0000000000000001",
48843 => "0000000000000001",48844 => "0000000000000001",
48845 => "0000000000000001",48846 => "0000000000000001",
48847 => "0000000000000001",48848 => "0000000000000001",
48849 => "0000000000000001",48850 => "0000000000000001",
48851 => "0000000000000001",48852 => "0000000000000001",
48853 => "0000000000000001",48854 => "0000000000000001",
48855 => "0000000000000001",48856 => "0000000000000001",
48857 => "0000000000000001",48858 => "0000000000000001",
48859 => "0000000000000001",48860 => "0000000000000001",
48861 => "0000000000000001",48862 => "0000000000000001",
48863 => "0000000000000001",48864 => "0000000000000001",
48865 => "0000000000000001",48866 => "0000000000000001",
48867 => "0000000000000001",48868 => "0000000000000001",
48869 => "0000000000000001",48870 => "0000000000000001",
48871 => "0000000000000001",48872 => "0000000000000001",
48873 => "0000000000000001",48874 => "0000000000000001",
48875 => "0000000000000001",48876 => "0000000000000001",
48877 => "0000000000000001",48878 => "0000000000000001",
48879 => "0000000000000001",48880 => "0000000000000001",
48881 => "0000000000000001",48882 => "0000000000000001",
48883 => "0000000000000001",48884 => "0000000000000001",
48885 => "0000000000000001",48886 => "0000000000000001",
48887 => "0000000000000001",48888 => "0000000000000001",
48889 => "0000000000000001",48890 => "0000000000000001",
48891 => "0000000000000001",48892 => "0000000000000001",
48893 => "0000000000000001",48894 => "0000000000000001",
48895 => "0000000000000001",48896 => "0000000000000001",
48897 => "0000000000000001",48898 => "0000000000000001",
48899 => "0000000000000001",48900 => "0000000000000001",
48901 => "0000000000000001",48902 => "0000000000000001",
48903 => "0000000000000001",48904 => "0000000000000001",
48905 => "0000000000000001",48906 => "0000000000000001",
48907 => "0000000000000001",48908 => "0000000000000001",
48909 => "0000000000000001",48910 => "0000000000000001",
48911 => "0000000000000001",48912 => "0000000000000001",
48913 => "0000000000000001",48914 => "0000000000000001",
48915 => "0000000000000001",48916 => "0000000000000001",
48917 => "0000000000000001",48918 => "0000000000000001",
48919 => "0000000000000001",48920 => "0000000000000001",
48921 => "0000000000000001",48922 => "0000000000000001",
48923 => "0000000000000001",48924 => "0000000000000001",
48925 => "0000000000000001",48926 => "0000000000000001",
48927 => "0000000000000001",48928 => "0000000000000001",
48929 => "0000000000000001",48930 => "0000000000000001",
48931 => "0000000000000001",48932 => "0000000000000001",
48933 => "0000000000000001",48934 => "0000000000000001",
48935 => "0000000000000001",48936 => "0000000000000001",
48937 => "0000000000000001",48938 => "0000000000000001",
48939 => "0000000000000001",48940 => "0000000000000001",
48941 => "0000000000000001",48942 => "0000000000000001",
48943 => "0000000000000001",48944 => "0000000000000001",
48945 => "0000000000000001",48946 => "0000000000000001",
48947 => "0000000000000001",48948 => "0000000000000001",
48949 => "0000000000000001",48950 => "0000000000000001",
48951 => "0000000000000001",48952 => "0000000000000001",
48953 => "0000000000000001",48954 => "0000000000000001",
48955 => "0000000000000001",48956 => "0000000000000001",
48957 => "0000000000000001",48958 => "0000000000000001",
48959 => "0000000000000001",48960 => "0000000000000001",
48961 => "0000000000000001",48962 => "0000000000000001",
48963 => "0000000000000001",48964 => "0000000000000001",
48965 => "0000000000000001",48966 => "0000000000000001",
48967 => "0000000000000001",48968 => "0000000000000001",
48969 => "0000000000000001",48970 => "0000000000000001",
48971 => "0000000000000001",48972 => "0000000000000001",
48973 => "0000000000000001",48974 => "0000000000000001",
48975 => "0000000000000001",48976 => "0000000000000001",
48977 => "0000000000000001",48978 => "0000000000000001",
48979 => "0000000000000001",48980 => "0000000000000001",
48981 => "0000000000000001",48982 => "0000000000000001",
48983 => "0000000000000001",48984 => "0000000000000001",
48985 => "0000000000000001",48986 => "0000000000000001",
48987 => "0000000000000001",48988 => "0000000000000001",
48989 => "0000000000000001",48990 => "0000000000000001",
48991 => "0000000000000001",48992 => "0000000000000001",
48993 => "0000000000000001",48994 => "0000000000000001",
48995 => "0000000000000001",48996 => "0000000000000001",
48997 => "0000000000000001",48998 => "0000000000000001",
48999 => "0000000000000001",49000 => "0000000000000001",
49001 => "0000000000000001",49002 => "0000000000000001",
49003 => "0000000000000001",49004 => "0000000000000001",
49005 => "0000000000000001",49006 => "0000000000000001",
49007 => "0000000000000001",49008 => "0000000000000001",
49009 => "0000000000000001",49010 => "0000000000000001",
49011 => "0000000000000001",49012 => "0000000000000001",
49013 => "0000000000000001",49014 => "0000000000000001",
49015 => "0000000000000001",49016 => "0000000000000001",
49017 => "0000000000000001",49018 => "0000000000000001",
49019 => "0000000000000001",49020 => "0000000000000001",
49021 => "0000000000000001",49022 => "0000000000000001",
49023 => "0000000000000001",49024 => "0000000000000001",
49025 => "0000000000000001",49026 => "0000000000000001",
49027 => "0000000000000001",49028 => "0000000000000001",
49029 => "0000000000000001",49030 => "0000000000000001",
49031 => "0000000000000001",49032 => "0000000000000001",
49033 => "0000000000000001",49034 => "0000000000000001",
49035 => "0000000000000001",49036 => "0000000000000001",
49037 => "0000000000000001",49038 => "0000000000000001",
49039 => "0000000000000001",49040 => "0000000000000001",
49041 => "0000000000000001",49042 => "0000000000000001",
49043 => "0000000000000001",49044 => "0000000000000001",
49045 => "0000000000000001",49046 => "0000000000000001",
49047 => "0000000000000001",49048 => "0000000000000001",
49049 => "0000000000000001",49050 => "0000000000000001",
49051 => "0000000000000001",49052 => "0000000000000001",
49053 => "0000000000000001",49054 => "0000000000000001",
49055 => "0000000000000001",49056 => "0000000000000001",
49057 => "0000000000000001",49058 => "0000000000000001",
49059 => "0000000000000001",49060 => "0000000000000001",
49061 => "0000000000000001",49062 => "0000000000000001",
49063 => "0000000000000001",49064 => "0000000000000001",
49065 => "0000000000000001",49066 => "0000000000000001",
49067 => "0000000000000001",49068 => "0000000000000001",
49069 => "0000000000000001",49070 => "0000000000000001",
49071 => "0000000000000001",49072 => "0000000000000001",
49073 => "0000000000000001",49074 => "0000000000000001",
49075 => "0000000000000001",49076 => "0000000000000001",
49077 => "0000000000000001",49078 => "0000000000000001",
49079 => "0000000000000001",49080 => "0000000000000001",
49081 => "0000000000000001",49082 => "0000000000000001",
49083 => "0000000000000001",49084 => "0000000000000001",
49085 => "0000000000000001",49086 => "0000000000000001",
49087 => "0000000000000001",49088 => "0000000000000001",
49089 => "0000000000000001",49090 => "0000000000000001",
49091 => "0000000000000001",49092 => "0000000000000001",
49093 => "0000000000000001",49094 => "0000000000000001",
49095 => "0000000000000001",49096 => "0000000000000001",
49097 => "0000000000000001",49098 => "0000000000000001",
49099 => "0000000000000001",49100 => "0000000000000001",
49101 => "0000000000000001",49102 => "0000000000000001",
49103 => "0000000000000001",49104 => "0000000000000001",
49105 => "0000000000000001",49106 => "0000000000000001",
49107 => "0000000000000001",49108 => "0000000000000001",
49109 => "0000000000000001",49110 => "0000000000000001",
49111 => "0000000000000001",49112 => "0000000000000001",
49113 => "0000000000000001",49114 => "0000000000000001",
49115 => "0000000000000001",49116 => "0000000000000001",
49117 => "0000000000000001",49118 => "0000000000000001",
49119 => "0000000000000001",49120 => "0000000000000001",
49121 => "0000000000000001",49122 => "0000000000000001",
49123 => "0000000000000001",49124 => "0000000000000001",
49125 => "0000000000000001",49126 => "0000000000000001",
49127 => "0000000000000001",49128 => "0000000000000001",
49129 => "0000000000000001",49130 => "0000000000000001",
49131 => "0000000000000001",49132 => "0000000000000001",
49133 => "0000000000000001",49134 => "0000000000000001",
49135 => "0000000000000001",49136 => "0000000000000001",
49137 => "0000000000000001",49138 => "0000000000000001",
49139 => "0000000000000001",49140 => "0000000000000001",
49141 => "0000000000000001",49142 => "0000000000000001",
49143 => "0000000000000001",49144 => "0000000000000001",
49145 => "0000000000000001",49146 => "0000000000000001",
49147 => "0000000000000001",49148 => "0000000000000001",
49149 => "0000000000000001",49150 => "0000000000000001",
49151 => "0000000000000001",49152 => "0000000000000000",
49153 => "0000000000000000",49154 => "0000000000000000",
49155 => "0000000000000000",49156 => "0000000000000000",
49157 => "0000000000000000",49158 => "0000000000000000",
49159 => "0000000000000000",49160 => "0000000000000000",
49161 => "0000000000000000",49162 => "0000000000000000",
49163 => "0000000000000000",49164 => "0000000000000000",
49165 => "0000000000000000",49166 => "0000000000000000",
49167 => "0000000000000000",49168 => "0000000000000000",
49169 => "0000000000000000",49170 => "0000000000000000",
49171 => "0000000000000000",49172 => "0000000000000000",
49173 => "0000000000000000",49174 => "0000000000000000",
49175 => "0000000000000000",49176 => "0000000000000000",
49177 => "0000000000000000",49178 => "0000000000000000",
49179 => "0000000000000000",49180 => "0000000000000000",
49181 => "0000000000000000",49182 => "0000000000000000",
49183 => "0000000000000000",49184 => "0000000000000000",
49185 => "0000000000000000",49186 => "0000000000000000",
49187 => "0000000000000000",49188 => "0000000000000000",
49189 => "0000000000000000",49190 => "0000000000000000",
49191 => "0000000000000000",49192 => "0000000000000000",
49193 => "0000000000000000",49194 => "0000000000000000",
49195 => "0000000000000000",49196 => "0000000000000000",
49197 => "0000000000000000",49198 => "0000000000000000",
49199 => "0000000000000000",49200 => "0000000000000000",
49201 => "0000000000000000",49202 => "0000000000000000",
49203 => "0000000000000000",49204 => "0000000000000000",
49205 => "0000000000000000",49206 => "0000000000000000",
49207 => "0000000000000000",49208 => "0000000000000000",
49209 => "0000000000000000",49210 => "0000000000000000",
49211 => "0000000000000000",49212 => "0000000000000000",
49213 => "0000000000000000",49214 => "0000000000000000",
49215 => "0000000000000000",49216 => "0000000000000000",
49217 => "0000000000000000",49218 => "0000000000000000",
49219 => "0000000000000000",49220 => "0000000000000000",
49221 => "0000000000000000",49222 => "0000000000000000",
49223 => "0000000000000000",49224 => "0000000000000000",
49225 => "0000000000000000",49226 => "0000000000000000",
49227 => "0000000000000000",49228 => "0000000000000000",
49229 => "0000000000000000",49230 => "0000000000000000",
49231 => "0000000000000000",49232 => "0000000000000000",
49233 => "0000000000000000",49234 => "0000000000000000",
49235 => "0000000000000000",49236 => "0000000000000000",
49237 => "0000000000000000",49238 => "0000000000000000",
49239 => "0000000000000000",49240 => "0000000000000000",
49241 => "0000000000000000",49242 => "0000000000000000",
49243 => "0000000000000000",49244 => "0000000000000000",
49245 => "0000000000000000",49246 => "0000000000000000",
49247 => "0000000000000000",49248 => "0000000000000000",
49249 => "0000000000000000",49250 => "0000000000000000",
49251 => "0000000000000000",49252 => "0000000000000000",
49253 => "0000000000000000",49254 => "0000000000000000",
49255 => "0000000000000000",49256 => "0000000000000000",
49257 => "0000000000000000",49258 => "0000000000000000",
49259 => "0000000000000000",49260 => "0000000000000000",
49261 => "0000000000000000",49262 => "0000000000000000",
49263 => "0000000000000000",49264 => "0000000000000000",
49265 => "0000000000000000",49266 => "0000000000000000",
49267 => "0000000000000000",49268 => "0000000000000000",
49269 => "0000000000000000",49270 => "0000000000000000",
49271 => "0000000000000000",49272 => "0000000000000000",
49273 => "0000000000000000",49274 => "0000000000000000",
49275 => "0000000000000000",49276 => "0000000000000000",
49277 => "0000000000000000",49278 => "0000000000000000",
49279 => "0000000000000000",49280 => "0000000000000000",
49281 => "0000000000000000",49282 => "0000000000000000",
49283 => "0000000000000000",49284 => "0000000000000000",
49285 => "0000000000000000",49286 => "0000000000000000",
49287 => "0000000000000000",49288 => "0000000000000000",
49289 => "0000000000000000",49290 => "0000000000000000",
49291 => "0000000000000000",49292 => "0000000000000000",
49293 => "0000000000000000",49294 => "0000000000000000",
49295 => "0000000000000000",49296 => "0000000000000000",
49297 => "0000000000000000",49298 => "0000000000000000",
49299 => "0000000000000000",49300 => "0000000000000000",
49301 => "0000000000000000",49302 => "0000000000000000",
49303 => "0000000000000000",49304 => "0000000000000000",
49305 => "0000000000000000",49306 => "0000000000000000",
49307 => "0000000000000000",49308 => "0000000000000000",
49309 => "0000000000000000",49310 => "0000000000000000",
49311 => "0000000000000000",49312 => "0000000000000000",
49313 => "0000000000000000",49314 => "0000000000000000",
49315 => "0000000000000000",49316 => "0000000000000000",
49317 => "0000000000000000",49318 => "0000000000000000",
49319 => "0000000000000000",49320 => "0000000000000000",
49321 => "0000000000000000",49322 => "0000000000000000",
49323 => "0000000000000000",49324 => "0000000000000000",
49325 => "0000000000000000",49326 => "0000000000000000",
49327 => "0000000000000000",49328 => "0000000000000000",
49329 => "0000000000000000",49330 => "0000000000000000",
49331 => "0000000000000000",49332 => "0000000000000000",
49333 => "0000000000000000",49334 => "0000000000000000",
49335 => "0000000000000000",49336 => "0000000000000000",
49337 => "0000000000000000",49338 => "0000000000000000",
49339 => "0000000000000000",49340 => "0000000000000000",
49341 => "0000000000000000",49342 => "0000000000000000",
49343 => "0000000000000000",49344 => "0000000000000000",
49345 => "0000000000000000",49346 => "0000000000000000",
49347 => "0000000000000000",49348 => "0000000000000000",
49349 => "0000000000000000",49350 => "0000000000000000",
49351 => "0000000000000000",49352 => "0000000000000000",
49353 => "0000000000000000",49354 => "0000000000000000",
49355 => "0000000000000000",49356 => "0000000000000000",
49357 => "0000000000000000",49358 => "0000000000000000",
49359 => "0000000000000000",49360 => "0000000000000000",
49361 => "0000000000000000",49362 => "0000000000000000",
49363 => "0000000000000000",49364 => "0000000000000000",
49365 => "0000000000000000",49366 => "0000000000000000",
49367 => "0000000000000000",49368 => "0000000000000000",
49369 => "0000000000000000",49370 => "0000000000000000",
49371 => "0000000000000000",49372 => "0000000000000000",
49373 => "0000000000000000",49374 => "0000000000000000",
49375 => "0000000000000000",49376 => "0000000000000000",
49377 => "0000000000000000",49378 => "0000000000000000",
49379 => "0000000000000000",49380 => "0000000000000000",
49381 => "0000000000000000",49382 => "0000000000000000",
49383 => "0000000000000000",49384 => "0000000000000000",
49385 => "0000000000000000",49386 => "0000000000000000",
49387 => "0000000000000000",49388 => "0000000000000000",
49389 => "0000000000000000",49390 => "0000000000000000",
49391 => "0000000000000000",49392 => "0000000000000000",
49393 => "0000000000000000",49394 => "0000000000000000",
49395 => "0000000000000000",49396 => "0000000000000000",
49397 => "0000000000000000",49398 => "0000000000000000",
49399 => "0000000000000000",49400 => "0000000000000000",
49401 => "0000000000000000",49402 => "0000000000000000",
49403 => "0000000000000000",49404 => "0000000000000000",
49405 => "0000000000000000",49406 => "0000000000000000",
49407 => "0000000000000000",49408 => "0000000000000000",
49409 => "0000000000000000",49410 => "0000000000000000",
49411 => "0000000000000000",49412 => "0000000000000000",
49413 => "0000000000000000",49414 => "0000000000000000",
49415 => "0000000000000000",49416 => "0000000000000000",
49417 => "0000000000000000",49418 => "0000000000000000",
49419 => "0000000000000000",49420 => "0000000000000000",
49421 => "0000000000000000",49422 => "0000000000000000",
49423 => "0000000000000000",49424 => "0000000000000000",
49425 => "0000000000000000",49426 => "0000000000000000",
49427 => "0000000000000000",49428 => "0000000000000000",
49429 => "0000000000000000",49430 => "0000000000000000",
49431 => "0000000000000000",49432 => "0000000000000000",
49433 => "0000000000000000",49434 => "0000000000000000",
49435 => "0000000000000000",49436 => "0000000000000000",
49437 => "0000000000000000",49438 => "0000000000000000",
49439 => "0000000000000000",49440 => "0000000000000000",
49441 => "0000000000000000",49442 => "0000000000000000",
49443 => "0000000000000000",49444 => "0000000000000000",
49445 => "0000000000000000",49446 => "0000000000000000",
49447 => "0000000000000000",49448 => "0000000000000000",
49449 => "0000000000000000",49450 => "0000000000000000",
49451 => "0000000000000000",49452 => "0000000000000000",
49453 => "0000000000000000",49454 => "0000000000000000",
49455 => "0000000000000000",49456 => "0000000000000000",
49457 => "0000000000000000",49458 => "0000000000000000",
49459 => "0000000000000000",49460 => "0000000000000000",
49461 => "0000000000000000",49462 => "0000000000000000",
49463 => "0000000000000000",49464 => "0000000000000000",
49465 => "0000000000000000",49466 => "0000000000000000",
49467 => "0000000000000000",49468 => "0000000000000000",
49469 => "0000000000000000",49470 => "0000000000000000",
49471 => "0000000000000000",49472 => "0000000000000000",
49473 => "0000000000000000",49474 => "0000000000000000",
49475 => "0000000000000000",49476 => "0000000000000000",
49477 => "0000000000000000",49478 => "0000000000000000",
49479 => "0000000000000000",49480 => "0000000000000000",
49481 => "0000000000000000",49482 => "0000000000000000",
49483 => "0000000000000000",49484 => "0000000000000000",
49485 => "0000000000000000",49486 => "0000000000000000",
49487 => "0000000000000000",49488 => "0000000000000000",
49489 => "0000000000000000",49490 => "0000000000000000",
49491 => "0000000000000000",49492 => "0000000000000000",
49493 => "0000000000000000",49494 => "0000000000000000",
49495 => "0000000000000000",49496 => "0000000000000000",
49497 => "0000000000000000",49498 => "0000000000000000",
49499 => "0000000000000000",49500 => "0000000000000000",
49501 => "0000000000000000",49502 => "0000000000000000",
49503 => "0000000000000000",49504 => "0000000000000000",
49505 => "0000000000000000",49506 => "0000000000000000",
49507 => "0000000000000000",49508 => "0000000000000000",
49509 => "0000000000000000",49510 => "0000000000000000",
49511 => "0000000000000000",49512 => "0000000000000000",
49513 => "0000000000000000",49514 => "0000000000000000",
49515 => "0000000000000000",49516 => "0000000000000000",
49517 => "0000000000000000",49518 => "0000000000000000",
49519 => "0000000000000000",49520 => "0000000000000000",
49521 => "0000000000000000",49522 => "0000000000000000",
49523 => "0000000000000000",49524 => "0000000000000000",
49525 => "0000000000000000",49526 => "0000000000000000",
49527 => "0000000000000000",49528 => "0000000000000000",
49529 => "0000000000000000",49530 => "0000000000000000",
49531 => "0000000000000000",49532 => "0000000000000000",
49533 => "0000000000000000",49534 => "0000000000000000",
49535 => "0000000000000000",49536 => "0000000000000000",
49537 => "0000000000000000",49538 => "0000000000000000",
49539 => "0000000000000000",49540 => "0000000000000000",
49541 => "0000000000000000",49542 => "0000000000000000",
49543 => "0000000000000000",49544 => "0000000000000000",
49545 => "0000000000000000",49546 => "0000000000000000",
49547 => "0000000000000000",49548 => "0000000000000000",
49549 => "0000000000000000",49550 => "0000000000000000",
49551 => "0000000000000000",49552 => "0000000000000000",
49553 => "0000000000000000",49554 => "0000000000000000",
49555 => "0000000000000000",49556 => "0000000000000000",
49557 => "0000000000000000",49558 => "0000000000000000",
49559 => "0000000000000000",49560 => "0000000000000000",
49561 => "0000000000000000",49562 => "0000000000000000",
49563 => "0000000000000000",49564 => "0000000000000000",
49565 => "0000000000000000",49566 => "0000000000000000",
49567 => "0000000000000000",49568 => "0000000000000000",
49569 => "0000000000000000",49570 => "0000000000000000",
49571 => "0000000000000000",49572 => "0000000000000000",
49573 => "0000000000000000",49574 => "0000000000000000",
49575 => "0000000000000000",49576 => "0000000000000000",
49577 => "0000000000000000",49578 => "0000000000000000",
49579 => "0000000000000000",49580 => "0000000000000000",
49581 => "0000000000000000",49582 => "0000000000000000",
49583 => "0000000000000000",49584 => "0000000000000000",
49585 => "0000000000000000",49586 => "0000000000000000",
49587 => "0000000000000000",49588 => "0000000000000000",
49589 => "0000000000000000",49590 => "0000000000000000",
49591 => "0000000000000000",49592 => "0000000000000000",
49593 => "0000000000000000",49594 => "0000000000000000",
49595 => "0000000000000000",49596 => "0000000000000000",
49597 => "0000000000000000",49598 => "0000000000000000",
49599 => "0000000000000000",49600 => "0000000000000000",
49601 => "0000000000000000",49602 => "0000000000000000",
49603 => "0000000000000000",49604 => "0000000000000000",
49605 => "0000000000000000",49606 => "0000000000000000",
49607 => "0000000000000000",49608 => "0000000000000000",
49609 => "0000000000000000",49610 => "0000000000000000",
49611 => "0000000000000000",49612 => "0000000000000000",
49613 => "0000000000000000",49614 => "0000000000000000",
49615 => "0000000000000000",49616 => "0000000000000000",
49617 => "0000000000000000",49618 => "0000000000000000",
49619 => "0000000000000000",49620 => "0000000000000000",
49621 => "0000000000000000",49622 => "0000000000000000",
49623 => "0000000000000000",49624 => "0000000000000000",
49625 => "0000000000000000",49626 => "0000000000000000",
49627 => "0000000000000000",49628 => "0000000000000000",
49629 => "0000000000000000",49630 => "0000000000000000",
49631 => "0000000000000000",49632 => "0000000000000000",
49633 => "0000000000000000",49634 => "0000000000000000",
49635 => "0000000000000000",49636 => "0000000000000000",
49637 => "0000000000000000",49638 => "0000000000000000",
49639 => "0000000000000000",49640 => "0000000000000000",
49641 => "0000000000000000",49642 => "0000000000000000",
49643 => "0000000000000000",49644 => "0000000000000000",
49645 => "0000000000000000",49646 => "0000000000000000",
49647 => "0000000000000000",49648 => "0000000000000000",
49649 => "0000000000000000",49650 => "0000000000000000",
49651 => "0000000000000000",49652 => "0000000000000000",
49653 => "0000000000000000",49654 => "0000000000000000",
49655 => "0000000000000000",49656 => "0000000000000000",
49657 => "0000000000000000",49658 => "0000000000000000",
49659 => "0000000000000000",49660 => "0000000000000000",
49661 => "0000000000000000",49662 => "0000000000000000",
49663 => "0000000000000000",49664 => "0000000000000000",
49665 => "0000000000000000",49666 => "0000000000000000",
49667 => "0000000000000000",49668 => "0000000000000000",
49669 => "0000000000000000",49670 => "0000000000000000",
49671 => "0000000000000000",49672 => "0000000000000000",
49673 => "0000000000000000",49674 => "0000000000000000",
49675 => "0000000000000000",49676 => "0000000000000000",
49677 => "0000000000000000",49678 => "0000000000000000",
49679 => "0000000000000000",49680 => "0000000000000000",
49681 => "0000000000000000",49682 => "0000000000000000",
49683 => "0000000000000000",49684 => "0000000000000000",
49685 => "0000000000000000",49686 => "0000000000000000",
49687 => "0000000000000000",49688 => "0000000000000000",
49689 => "0000000000000000",49690 => "0000000000000000",
49691 => "0000000000000000",49692 => "0000000000000000",
49693 => "0000000000000000",49694 => "0000000000000000",
49695 => "0000000000000000",49696 => "0000000000000000",
49697 => "0000000000000000",49698 => "0000000000000000",
49699 => "0000000000000000",49700 => "0000000000000000",
49701 => "0000000000000000",49702 => "0000000000000000",
49703 => "0000000000000000",49704 => "0000000000000000",
49705 => "0000000000000000",49706 => "0000000000000000",
49707 => "0000000000000000",49708 => "0000000000000000",
49709 => "0000000000000000",49710 => "0000000000000000",
49711 => "0000000000000000",49712 => "0000000000000000",
49713 => "0000000000000000",49714 => "0000000000000000",
49715 => "0000000000000000",49716 => "0000000000000000",
49717 => "0000000000000000",49718 => "0000000000000000",
49719 => "0000000000000000",49720 => "0000000000000000",
49721 => "0000000000000000",49722 => "0000000000000000",
49723 => "0000000000000000",49724 => "0000000000000000",
49725 => "0000000000000000",49726 => "0000000000000000",
49727 => "0000000000000000",49728 => "0000000000000000",
49729 => "0000000000000000",49730 => "0000000000000000",
49731 => "0000000000000000",49732 => "0000000000000000",
49733 => "0000000000000000",49734 => "0000000000000000",
49735 => "0000000000000000",49736 => "0000000000000000",
49737 => "0000000000000000",49738 => "0000000000000000",
49739 => "0000000000000000",49740 => "0000000000000000",
49741 => "0000000000000000",49742 => "0000000000000000",
49743 => "0000000000000000",49744 => "0000000000000000",
49745 => "0000000000000000",49746 => "0000000000000000",
49747 => "0000000000000000",49748 => "0000000000000000",
49749 => "0000000000000000",49750 => "0000000000000000",
49751 => "0000000000000000",49752 => "0000000000000000",
49753 => "0000000000000000",49754 => "0000000000000000",
49755 => "0000000000000000",49756 => "0000000000000000",
49757 => "0000000000000000",49758 => "0000000000000000",
49759 => "0000000000000000",49760 => "0000000000000000",
49761 => "0000000000000000",49762 => "0000000000000000",
49763 => "0000000000000000",49764 => "0000000000000000",
49765 => "0000000000000000",49766 => "0000000000000000",
49767 => "0000000000000000",49768 => "0000000000000000",
49769 => "0000000000000000",49770 => "0000000000000000",
49771 => "0000000000000000",49772 => "0000000000000000",
49773 => "0000000000000000",49774 => "0000000000000000",
49775 => "0000000000000000",49776 => "0000000000000000",
49777 => "0000000000000000",49778 => "0000000000000000",
49779 => "0000000000000000",49780 => "0000000000000000",
49781 => "0000000000000000",49782 => "0000000000000000",
49783 => "0000000000000000",49784 => "0000000000000000",
49785 => "0000000000000000",49786 => "0000000000000000",
49787 => "0000000000000000",49788 => "0000000000000000",
49789 => "0000000000000000",49790 => "0000000000000000",
49791 => "0000000000000000",49792 => "0000000000000000",
49793 => "0000000000000000",49794 => "0000000000000000",
49795 => "0000000000000000",49796 => "0000000000000000",
49797 => "0000000000000000",49798 => "0000000000000000",
49799 => "0000000000000000",49800 => "0000000000000000",
49801 => "0000000000000000",49802 => "0000000000000000",
49803 => "0000000000000000",49804 => "0000000000000000",
49805 => "0000000000000000",49806 => "0000000000000000",
49807 => "0000000000000000",49808 => "0000000000000000",
49809 => "0000000000000000",49810 => "0000000000000000",
49811 => "0000000000000000",49812 => "0000000000000000",
49813 => "0000000000000000",49814 => "0000000000000000",
49815 => "0000000000000000",49816 => "0000000000000000",
49817 => "0000000000000000",49818 => "0000000000000000",
49819 => "0000000000000000",49820 => "0000000000000000",
49821 => "0000000000000000",49822 => "0000000000000000",
49823 => "0000000000000000",49824 => "0000000000000000",
49825 => "0000000000000000",49826 => "0000000000000000",
49827 => "0000000000000000",49828 => "0000000000000000",
49829 => "0000000000000000",49830 => "0000000000000000",
49831 => "0000000000000000",49832 => "0000000000000000",
49833 => "0000000000000000",49834 => "0000000000000000",
49835 => "0000000000000000",49836 => "0000000000000000",
49837 => "0000000000000000",49838 => "0000000000000000",
49839 => "0000000000000000",49840 => "0000000000000000",
49841 => "0000000000000000",49842 => "0000000000000000",
49843 => "0000000000000000",49844 => "0000000000000000",
49845 => "0000000000000000",49846 => "0000000000000000",
49847 => "0000000000000000",49848 => "0000000000000000",
49849 => "0000000000000000",49850 => "0000000000000000",
49851 => "0000000000000000",49852 => "0000000000000000",
49853 => "0000000000000000",49854 => "0000000000000000",
49855 => "0000000000000000",49856 => "0000000000000000",
49857 => "0000000000000000",49858 => "0000000000000000",
49859 => "0000000000000000",49860 => "0000000000000000",
49861 => "0000000000000000",49862 => "0000000000000000",
49863 => "0000000000000000",49864 => "0000000000000000",
49865 => "0000000000000000",49866 => "0000000000000000",
49867 => "0000000000000000",49868 => "0000000000000000",
49869 => "0000000000000000",49870 => "0000000000000000",
49871 => "0000000000000000",49872 => "0000000000000000",
49873 => "0000000000000000",49874 => "0000000000000000",
49875 => "0000000000000000",49876 => "0000000000000000",
49877 => "0000000000000000",49878 => "0000000000000000",
49879 => "0000000000000000",49880 => "0000000000000000",
49881 => "0000000000000000",49882 => "0000000000000000",
49883 => "0000000000000000",49884 => "0000000000000000",
49885 => "0000000000000000",49886 => "0000000000000000",
49887 => "0000000000000000",49888 => "0000000000000000",
49889 => "0000000000000000",49890 => "0000000000000000",
49891 => "0000000000000000",49892 => "0000000000000000",
49893 => "0000000000000000",49894 => "0000000000000000",
49895 => "0000000000000000",49896 => "0000000000000000",
49897 => "0000000000000000",49898 => "0000000000000000",
49899 => "0000000000000000",49900 => "0000000000000000",
49901 => "0000000000000000",49902 => "0000000000000000",
49903 => "0000000000000000",49904 => "0000000000000000",
49905 => "0000000000000000",49906 => "0000000000000000",
49907 => "0000000000000000",49908 => "0000000000000000",
49909 => "0000000000000000",49910 => "0000000000000000",
49911 => "0000000000000000",49912 => "0000000000000000",
49913 => "0000000000000000",49914 => "0000000000000000",
49915 => "0000000000000000",49916 => "0000000000000000",
49917 => "0000000000000000",49918 => "0000000000000000",
49919 => "0000000000000000",49920 => "0000000000000000",
49921 => "0000000000000000",49922 => "0000000000000000",
49923 => "0000000000000000",49924 => "0000000000000000",
49925 => "0000000000000000",49926 => "0000000000000000",
49927 => "0000000000000000",49928 => "0000000000000000",
49929 => "0000000000000000",49930 => "0000000000000000",
49931 => "0000000000000000",49932 => "0000000000000000",
49933 => "0000000000000000",49934 => "0000000000000000",
49935 => "0000000000000000",49936 => "0000000000000000",
49937 => "0000000000000000",49938 => "0000000000000000",
49939 => "0000000000000000",49940 => "0000000000000000",
49941 => "0000000000000000",49942 => "0000000000000000",
49943 => "0000000000000000",49944 => "0000000000000000",
49945 => "0000000000000000",49946 => "0000000000000000",
49947 => "0000000000000000",49948 => "0000000000000000",
49949 => "0000000000000000",49950 => "0000000000000000",
49951 => "0000000000000000",49952 => "0000000000000000",
49953 => "0000000000000000",49954 => "0000000000000000",
49955 => "0000000000000000",49956 => "0000000000000000",
49957 => "0000000000000000",49958 => "0000000000000000",
49959 => "0000000000000000",49960 => "0000000000000000",
49961 => "0000000000000000",49962 => "0000000000000000",
49963 => "0000000000000000",49964 => "0000000000000000",
49965 => "0000000000000000",49966 => "0000000000000000",
49967 => "0000000000000000",49968 => "0000000000000000",
49969 => "0000000000000000",49970 => "0000000000000000",
49971 => "0000000000000000",49972 => "0000000000000000",
49973 => "0000000000000000",49974 => "0000000000000000",
49975 => "0000000000000000",49976 => "0000000000000000",
49977 => "0000000000000000",49978 => "0000000000000000",
49979 => "0000000000000000",49980 => "0000000000000000",
49981 => "0000000000000000",49982 => "0000000000000000",
49983 => "0000000000000000",49984 => "0000000000000000",
49985 => "0000000000000000",49986 => "0000000000000000",
49987 => "0000000000000000",49988 => "0000000000000000",
49989 => "0000000000000000",49990 => "0000000000000000",
49991 => "0000000000000000",49992 => "0000000000000000",
49993 => "0000000000000000",49994 => "0000000000000000",
49995 => "0000000000000000",49996 => "0000000000000000",
49997 => "0000000000000000",49998 => "0000000000000000",
49999 => "0000000000000000",50000 => "0000000000000000",
50001 => "0000000000000000",50002 => "0000000000000000",
50003 => "0000000000000000",50004 => "0000000000000000",
50005 => "0000000000000000",50006 => "0000000000000000",
50007 => "0000000000000000",50008 => "0000000000000000",
50009 => "0000000000000000",50010 => "0000000000000000",
50011 => "0000000000000000",50012 => "0000000000000000",
50013 => "0000000000000000",50014 => "0000000000000000",
50015 => "0000000000000000",50016 => "0000000000000000",
50017 => "0000000000000000",50018 => "0000000000000000",
50019 => "0000000000000000",50020 => "0000000000000000",
50021 => "0000000000000000",50022 => "0000000000000000",
50023 => "0000000000000000",50024 => "0000000000000000",
50025 => "0000000000000000",50026 => "0000000000000000",
50027 => "0000000000000000",50028 => "0000000000000000",
50029 => "0000000000000000",50030 => "0000000000000000",
50031 => "0000000000000000",50032 => "0000000000000000",
50033 => "0000000000000000",50034 => "0000000000000000",
50035 => "0000000000000000",50036 => "0000000000000000",
50037 => "0000000000000000",50038 => "0000000000000000",
50039 => "0000000000000000",50040 => "0000000000000000",
50041 => "0000000000000000",50042 => "0000000000000000",
50043 => "0000000000000000",50044 => "0000000000000000",
50045 => "0000000000000000",50046 => "0000000000000000",
50047 => "0000000000000000",50048 => "0000000000000000",
50049 => "0000000000000000",50050 => "0000000000000000",
50051 => "0000000000000000",50052 => "0000000000000000",
50053 => "0000000000000000",50054 => "0000000000000000",
50055 => "0000000000000000",50056 => "0000000000000000",
50057 => "0000000000000000",50058 => "0000000000000000",
50059 => "0000000000000000",50060 => "0000000000000000",
50061 => "0000000000000000",50062 => "0000000000000000",
50063 => "0000000000000000",50064 => "0000000000000000",
50065 => "0000000000000000",50066 => "0000000000000000",
50067 => "0000000000000000",50068 => "0000000000000000",
50069 => "0000000000000000",50070 => "0000000000000000",
50071 => "0000000000000000",50072 => "0000000000000000",
50073 => "0000000000000000",50074 => "0000000000000000",
50075 => "0000000000000000",50076 => "0000000000000000",
50077 => "0000000000000000",50078 => "0000000000000000",
50079 => "0000000000000000",50080 => "0000000000000000",
50081 => "0000000000000000",50082 => "0000000000000000",
50083 => "0000000000000000",50084 => "0000000000000000",
50085 => "0000000000000000",50086 => "0000000000000000",
50087 => "0000000000000000",50088 => "0000000000000000",
50089 => "0000000000000000",50090 => "0000000000000000",
50091 => "0000000000000000",50092 => "0000000000000000",
50093 => "0000000000000000",50094 => "0000000000000000",
50095 => "0000000000000000",50096 => "0000000000000000",
50097 => "0000000000000000",50098 => "0000000000000000",
50099 => "0000000000000000",50100 => "0000000000000000",
50101 => "0000000000000000",50102 => "0000000000000000",
50103 => "0000000000000000",50104 => "0000000000000000",
50105 => "0000000000000000",50106 => "0000000000000000",
50107 => "0000000000000000",50108 => "0000000000000000",
50109 => "0000000000000000",50110 => "0000000000000000",
50111 => "0000000000000000",50112 => "0000000000000000",
50113 => "0000000000000000",50114 => "0000000000000000",
50115 => "0000000000000000",50116 => "0000000000000000",
50117 => "0000000000000000",50118 => "0000000000000000",
50119 => "0000000000000000",50120 => "0000000000000000",
50121 => "0000000000000000",50122 => "0000000000000000",
50123 => "0000000000000000",50124 => "0000000000000000",
50125 => "0000000000000000",50126 => "0000000000000000",
50127 => "0000000000000000",50128 => "0000000000000000",
50129 => "0000000000000000",50130 => "0000000000000000",
50131 => "0000000000000000",50132 => "0000000000000000",
50133 => "0000000000000000",50134 => "0000000000000000",
50135 => "0000000000000000",50136 => "0000000000000000",
50137 => "0000000000000000",50138 => "0000000000000000",
50139 => "0000000000000000",50140 => "0000000000000000",
50141 => "0000000000000000",50142 => "0000000000000000",
50143 => "0000000000000000",50144 => "0000000000000000",
50145 => "0000000000000000",50146 => "0000000000000000",
50147 => "0000000000000000",50148 => "0000000000000000",
50149 => "0000000000000000",50150 => "0000000000000000",
50151 => "0000000000000000",50152 => "0000000000000000",
50153 => "0000000000000000",50154 => "0000000000000000",
50155 => "0000000000000000",50156 => "0000000000000000",
50157 => "0000000000000000",50158 => "0000000000000000",
50159 => "0000000000000000",50160 => "0000000000000000",
50161 => "0000000000000000",50162 => "0000000000000000",
50163 => "0000000000000000",50164 => "0000000000000000",
50165 => "0000000000000000",50166 => "0000000000000000",
50167 => "0000000000000000",50168 => "0000000000000000",
50169 => "0000000000000000",50170 => "0000000000000000",
50171 => "0000000000000000",50172 => "0000000000000000",
50173 => "0000000000000000",50174 => "0000000000000000",
50175 => "0000000000000000",50176 => "0000000000000000",
50177 => "0000000000000000",50178 => "0000000000000000",
50179 => "0000000000000000",50180 => "0000000000000000",
50181 => "0000000000000000",50182 => "0000000000000000",
50183 => "0000000000000000",50184 => "0000000000000000",
50185 => "0000000000000000",50186 => "0000000000000000",
50187 => "0000000000000000",50188 => "0000000000000000",
50189 => "0000000000000000",50190 => "0000000000000000",
50191 => "0000000000000000",50192 => "0000000000000000",
50193 => "0000000000000000",50194 => "0000000000000000",
50195 => "0000000000000000",50196 => "0000000000000000",
50197 => "0000000000000000",50198 => "0000000000000000",
50199 => "0000000000000000",50200 => "0000000000000000",
50201 => "0000000000000000",50202 => "0000000000000000",
50203 => "0000000000000000",50204 => "0000000000000000",
50205 => "0000000000000000",50206 => "0000000000000000",
50207 => "0000000000000000",50208 => "0000000000000000",
50209 => "0000000000000000",50210 => "0000000000000000",
50211 => "0000000000000000",50212 => "0000000000000000",
50213 => "0000000000000000",50214 => "0000000000000000",
50215 => "0000000000000000",50216 => "0000000000000000",
50217 => "0000000000000000",50218 => "0000000000000000",
50219 => "0000000000000000",50220 => "0000000000000000",
50221 => "0000000000000000",50222 => "0000000000000000",
50223 => "0000000000000000",50224 => "0000000000000000",
50225 => "0000000000000000",50226 => "0000000000000000",
50227 => "0000000000000000",50228 => "0000000000000000",
50229 => "0000000000000000",50230 => "0000000000000000",
50231 => "0000000000000000",50232 => "0000000000000000",
50233 => "0000000000000000",50234 => "0000000000000000",
50235 => "0000000000000000",50236 => "0000000000000000",
50237 => "0000000000000000",50238 => "0000000000000000",
50239 => "0000000000000000",50240 => "0000000000000000",
50241 => "0000000000000000",50242 => "0000000000000000",
50243 => "0000000000000000",50244 => "0000000000000000",
50245 => "0000000000000000",50246 => "0000000000000000",
50247 => "0000000000000000",50248 => "0000000000000000",
50249 => "0000000000000000",50250 => "0000000000000000",
50251 => "0000000000000000",50252 => "0000000000000000",
50253 => "0000000000000000",50254 => "0000000000000000",
50255 => "0000000000000000",50256 => "0000000000000000",
50257 => "0000000000000000",50258 => "0000000000000000",
50259 => "0000000000000000",50260 => "0000000000000000",
50261 => "0000000000000000",50262 => "0000000000000000",
50263 => "0000000000000000",50264 => "0000000000000000",
50265 => "0000000000000000",50266 => "0000000000000000",
50267 => "0000000000000000",50268 => "0000000000000000",
50269 => "0000000000000000",50270 => "0000000000000000",
50271 => "0000000000000000",50272 => "0000000000000000",
50273 => "0000000000000000",50274 => "0000000000000000",
50275 => "0000000000000000",50276 => "0000000000000000",
50277 => "0000000000000000",50278 => "0000000000000000",
50279 => "0000000000000000",50280 => "0000000000000000",
50281 => "0000000000000000",50282 => "0000000000000000",
50283 => "0000000000000000",50284 => "0000000000000000",
50285 => "0000000000000000",50286 => "0000000000000000",
50287 => "0000000000000000",50288 => "0000000000000000",
50289 => "0000000000000000",50290 => "0000000000000000",
50291 => "0000000000000000",50292 => "0000000000000000",
50293 => "0000000000000000",50294 => "0000000000000000",
50295 => "0000000000000000",50296 => "0000000000000000",
50297 => "0000000000000000",50298 => "0000000000000000",
50299 => "0000000000000000",50300 => "0000000000000000",
50301 => "0000000000000000",50302 => "0000000000000000",
50303 => "0000000000000000",50304 => "0000000000000000",
50305 => "0000000000000000",50306 => "0000000000000000",
50307 => "0000000000000000",50308 => "0000000000000000",
50309 => "0000000000000000",50310 => "0000000000000000",
50311 => "0000000000000000",50312 => "0000000000000000",
50313 => "0000000000000000",50314 => "0000000000000000",
50315 => "0000000000000000",50316 => "0000000000000000",
50317 => "0000000000000000",50318 => "0000000000000000",
50319 => "0000000000000000",50320 => "0000000000000000",
50321 => "0000000000000000",50322 => "0000000000000000",
50323 => "0000000000000000",50324 => "0000000000000000",
50325 => "0000000000000000",50326 => "0000000000000000",
50327 => "0000000000000000",50328 => "0000000000000000",
50329 => "0000000000000000",50330 => "0000000000000000",
50331 => "0000000000000000",50332 => "0000000000000000",
50333 => "0000000000000000",50334 => "0000000000000000",
50335 => "0000000000000000",50336 => "0000000000000000",
50337 => "0000000000000000",50338 => "0000000000000000",
50339 => "0000000000000000",50340 => "0000000000000000",
50341 => "0000000000000000",50342 => "0000000000000000",
50343 => "0000000000000000",50344 => "0000000000000000",
50345 => "0000000000000000",50346 => "0000000000000000",
50347 => "0000000000000000",50348 => "0000000000000000",
50349 => "0000000000000000",50350 => "0000000000000000",
50351 => "0000000000000000",50352 => "0000000000000000",
50353 => "0000000000000000",50354 => "0000000000000000",
50355 => "0000000000000000",50356 => "0000000000000000",
50357 => "0000000000000000",50358 => "0000000000000000",
50359 => "0000000000000000",50360 => "0000000000000000",
50361 => "0000000000000000",50362 => "0000000000000000",
50363 => "0000000000000000",50364 => "0000000000000000",
50365 => "0000000000000000",50366 => "0000000000000000",
50367 => "0000000000000000",50368 => "0000000000000000",
50369 => "0000000000000000",50370 => "0000000000000000",
50371 => "0000000000000000",50372 => "0000000000000000",
50373 => "0000000000000000",50374 => "0000000000000000",
50375 => "0000000000000000",50376 => "0000000000000000",
50377 => "0000000000000000",50378 => "0000000000000000",
50379 => "0000000000000000",50380 => "0000000000000000",
50381 => "0000000000000000",50382 => "0000000000000000",
50383 => "0000000000000000",50384 => "0000000000000000",
50385 => "0000000000000000",50386 => "0000000000000000",
50387 => "0000000000000000",50388 => "0000000000000000",
50389 => "0000000000000000",50390 => "0000000000000000",
50391 => "0000000000000000",50392 => "0000000000000000",
50393 => "0000000000000000",50394 => "0000000000000000",
50395 => "0000000000000000",50396 => "0000000000000000",
50397 => "0000000000000000",50398 => "0000000000000000",
50399 => "0000000000000000",50400 => "0000000000000000",
50401 => "0000000000000000",50402 => "0000000000000000",
50403 => "0000000000000000",50404 => "0000000000000000",
50405 => "0000000000000000",50406 => "0000000000000000",
50407 => "0000000000000000",50408 => "0000000000000000",
50409 => "0000000000000000",50410 => "0000000000000000",
50411 => "0000000000000000",50412 => "0000000000000000",
50413 => "0000000000000000",50414 => "0000000000000000",
50415 => "0000000000000000",50416 => "0000000000000000",
50417 => "0000000000000000",50418 => "0000000000000000",
50419 => "0000000000000000",50420 => "0000000000000000",
50421 => "0000000000000000",50422 => "0000000000000000",
50423 => "0000000000000000",50424 => "0000000000000000",
50425 => "0000000000000000",50426 => "0000000000000000",
50427 => "0000000000000000",50428 => "0000000000000000",
50429 => "0000000000000000",50430 => "0000000000000000",
50431 => "0000000000000000",50432 => "0000000000000000",
50433 => "0000000000000000",50434 => "0000000000000000",
50435 => "0000000000000000",50436 => "0000000000000000",
50437 => "0000000000000000",50438 => "0000000000000000",
50439 => "0000000000000000",50440 => "0000000000000000",
50441 => "0000000000000000",50442 => "0000000000000000",
50443 => "0000000000000000",50444 => "0000000000000000",
50445 => "0000000000000000",50446 => "0000000000000000",
50447 => "0000000000000000",50448 => "0000000000000000",
50449 => "0000000000000000",50450 => "0000000000000000",
50451 => "0000000000000000",50452 => "0000000000000000",
50453 => "0000000000000000",50454 => "0000000000000000",
50455 => "0000000000000000",50456 => "0000000000000000",
50457 => "0000000000000000",50458 => "0000000000000000",
50459 => "0000000000000000",50460 => "0000000000000000",
50461 => "0000000000000000",50462 => "0000000000000000",
50463 => "0000000000000000",50464 => "0000000000000000",
50465 => "0000000000000000",50466 => "0000000000000000",
50467 => "0000000000000000",50468 => "0000000000000000",
50469 => "0000000000000000",50470 => "0000000000000000",
50471 => "0000000000000000",50472 => "0000000000000000",
50473 => "0000000000000000",50474 => "0000000000000000",
50475 => "0000000000000000",50476 => "0000000000000000",
50477 => "0000000000000000",50478 => "0000000000000000",
50479 => "0000000000000000",50480 => "0000000000000000",
50481 => "0000000000000000",50482 => "0000000000000000",
50483 => "0000000000000000",50484 => "0000000000000000",
50485 => "0000000000000000",50486 => "0000000000000000",
50487 => "0000000000000000",50488 => "0000000000000000",
50489 => "0000000000000000",50490 => "0000000000000000",
50491 => "0000000000000000",50492 => "0000000000000000",
50493 => "0000000000000000",50494 => "0000000000000000",
50495 => "0000000000000000",50496 => "0000000000000000",
50497 => "0000000000000000",50498 => "0000000000000000",
50499 => "0000000000000000",50500 => "0000000000000000",
50501 => "0000000000000000",50502 => "0000000000000000",
50503 => "0000000000000000",50504 => "0000000000000000",
50505 => "0000000000000000",50506 => "0000000000000000",
50507 => "0000000000000000",50508 => "0000000000000000",
50509 => "0000000000000000",50510 => "0000000000000000",
50511 => "0000000000000000",50512 => "0000000000000000",
50513 => "0000000000000000",50514 => "0000000000000000",
50515 => "0000000000000000",50516 => "0000000000000000",
50517 => "0000000000000000",50518 => "0000000000000000",
50519 => "0000000000000000",50520 => "0000000000000000",
50521 => "0000000000000000",50522 => "0000000000000000",
50523 => "0000000000000000",50524 => "0000000000000000",
50525 => "0000000000000000",50526 => "0000000000000000",
50527 => "0000000000000000",50528 => "0000000000000000",
50529 => "0000000000000000",50530 => "0000000000000000",
50531 => "0000000000000000",50532 => "0000000000000000",
50533 => "0000000000000000",50534 => "0000000000000000",
50535 => "0000000000000000",50536 => "0000000000000000",
50537 => "0000000000000000",50538 => "0000000000000000",
50539 => "0000000000000000",50540 => "0000000000000000",
50541 => "0000000000000000",50542 => "0000000000000000",
50543 => "0000000000000000",50544 => "0000000000000000",
50545 => "0000000000000000",50546 => "0000000000000000",
50547 => "0000000000000000",50548 => "0000000000000000",
50549 => "0000000000000000",50550 => "0000000000000000",
50551 => "0000000000000000",50552 => "0000000000000000",
50553 => "0000000000000000",50554 => "0000000000000000",
50555 => "0000000000000000",50556 => "0000000000000000",
50557 => "0000000000000000",50558 => "0000000000000000",
50559 => "0000000000000000",50560 => "0000000000000000",
50561 => "0000000000000000",50562 => "0000000000000000",
50563 => "0000000000000000",50564 => "0000000000000000",
50565 => "0000000000000000",50566 => "0000000000000000",
50567 => "0000000000000000",50568 => "0000000000000000",
50569 => "0000000000000000",50570 => "0000000000000000",
50571 => "0000000000000000",50572 => "0000000000000000",
50573 => "0000000000000000",50574 => "0000000000000000",
50575 => "0000000000000000",50576 => "0000000000000000",
50577 => "0000000000000000",50578 => "0000000000000000",
50579 => "0000000000000000",50580 => "0000000000000000",
50581 => "0000000000000000",50582 => "0000000000000000",
50583 => "0000000000000000",50584 => "0000000000000000",
50585 => "0000000000000000",50586 => "0000000000000000",
50587 => "0000000000000000",50588 => "0000000000000000",
50589 => "0000000000000000",50590 => "0000000000000000",
50591 => "0000000000000000",50592 => "0000000000000000",
50593 => "0000000000000000",50594 => "0000000000000000",
50595 => "0000000000000000",50596 => "0000000000000000",
50597 => "0000000000000000",50598 => "0000000000000000",
50599 => "0000000000000000",50600 => "0000000000000000",
50601 => "0000000000000000",50602 => "0000000000000000",
50603 => "0000000000000000",50604 => "0000000000000000",
50605 => "0000000000000000",50606 => "0000000000000000",
50607 => "0000000000000000",50608 => "0000000000000000",
50609 => "0000000000000000",50610 => "0000000000000000",
50611 => "0000000000000000",50612 => "0000000000000000",
50613 => "0000000000000000",50614 => "0000000000000000",
50615 => "0000000000000000",50616 => "0000000000000000",
50617 => "0000000000000000",50618 => "0000000000000000",
50619 => "0000000000000000",50620 => "0000000000000000",
50621 => "0000000000000000",50622 => "0000000000000000",
50623 => "0000000000000000",50624 => "0000000000000000",
50625 => "0000000000000000",50626 => "0000000000000000",
50627 => "0000000000000000",50628 => "0000000000000000",
50629 => "0000000000000000",50630 => "0000000000000000",
50631 => "0000000000000000",50632 => "0000000000000000",
50633 => "0000000000000000",50634 => "0000000000000000",
50635 => "0000000000000000",50636 => "0000000000000000",
50637 => "0000000000000000",50638 => "0000000000000000",
50639 => "0000000000000000",50640 => "0000000000000000",
50641 => "0000000000000000",50642 => "0000000000000000",
50643 => "0000000000000000",50644 => "0000000000000000",
50645 => "0000000000000000",50646 => "0000000000000000",
50647 => "0000000000000000",50648 => "0000000000000000",
50649 => "0000000000000000",50650 => "0000000000000000",
50651 => "0000000000000000",50652 => "0000000000000000",
50653 => "0000000000000000",50654 => "0000000000000000",
50655 => "0000000000000000",50656 => "0000000000000000",
50657 => "0000000000000000",50658 => "0000000000000000",
50659 => "0000000000000000",50660 => "0000000000000000",
50661 => "0000000000000000",50662 => "0000000000000000",
50663 => "0000000000000000",50664 => "0000000000000000",
50665 => "0000000000000000",50666 => "0000000000000000",
50667 => "0000000000000000",50668 => "0000000000000000",
50669 => "0000000000000000",50670 => "0000000000000000",
50671 => "0000000000000000",50672 => "0000000000000000",
50673 => "0000000000000000",50674 => "0000000000000000",
50675 => "0000000000000000",50676 => "0000000000000000",
50677 => "0000000000000000",50678 => "0000000000000000",
50679 => "0000000000000000",50680 => "0000000000000000",
50681 => "0000000000000000",50682 => "0000000000000000",
50683 => "0000000000000000",50684 => "0000000000000000",
50685 => "0000000000000000",50686 => "0000000000000000",
50687 => "0000000000000000",50688 => "0000000000000000",
50689 => "0000000000000000",50690 => "0000000000000000",
50691 => "0000000000000000",50692 => "0000000000000000",
50693 => "0000000000000000",50694 => "0000000000000000",
50695 => "0000000000000000",50696 => "0000000000000000",
50697 => "0000000000000000",50698 => "0000000000000000",
50699 => "0000000000000000",50700 => "0000000000000000",
50701 => "0000000000000000",50702 => "0000000000000000",
50703 => "0000000000000000",50704 => "0000000000000000",
50705 => "0000000000000000",50706 => "0000000000000000",
50707 => "0000000000000000",50708 => "0000000000000000",
50709 => "0000000000000000",50710 => "0000000000000000",
50711 => "0000000000000000",50712 => "0000000000000000",
50713 => "0000000000000000",50714 => "0000000000000000",
50715 => "0000000000000000",50716 => "0000000000000000",
50717 => "0000000000000000",50718 => "0000000000000000",
50719 => "0000000000000000",50720 => "0000000000000000",
50721 => "0000000000000000",50722 => "0000000000000000",
50723 => "0000000000000000",50724 => "0000000000000000",
50725 => "0000000000000000",50726 => "0000000000000000",
50727 => "0000000000000000",50728 => "0000000000000000",
50729 => "0000000000000000",50730 => "0000000000000000",
50731 => "0000000000000000",50732 => "0000000000000000",
50733 => "0000000000000000",50734 => "0000000000000000",
50735 => "0000000000000000",50736 => "0000000000000000",
50737 => "0000000000000000",50738 => "0000000000000000",
50739 => "0000000000000000",50740 => "0000000000000000",
50741 => "0000000000000000",50742 => "0000000000000000",
50743 => "0000000000000000",50744 => "0000000000000000",
50745 => "0000000000000000",50746 => "0000000000000000",
50747 => "0000000000000000",50748 => "0000000000000000",
50749 => "0000000000000000",50750 => "0000000000000000",
50751 => "0000000000000000",50752 => "0000000000000000",
50753 => "0000000000000000",50754 => "0000000000000000",
50755 => "0000000000000000",50756 => "0000000000000000",
50757 => "0000000000000000",50758 => "0000000000000000",
50759 => "0000000000000000",50760 => "0000000000000000",
50761 => "0000000000000000",50762 => "0000000000000000",
50763 => "0000000000000000",50764 => "0000000000000000",
50765 => "0000000000000000",50766 => "0000000000000000",
50767 => "0000000000000000",50768 => "0000000000000000",
50769 => "0000000000000000",50770 => "0000000000000000",
50771 => "0000000000000000",50772 => "0000000000000000",
50773 => "0000000000000000",50774 => "0000000000000000",
50775 => "0000000000000000",50776 => "0000000000000000",
50777 => "0000000000000000",50778 => "0000000000000000",
50779 => "0000000000000000",50780 => "0000000000000000",
50781 => "0000000000000000",50782 => "0000000000000000",
50783 => "0000000000000000",50784 => "0000000000000000",
50785 => "0000000000000000",50786 => "0000000000000000",
50787 => "0000000000000000",50788 => "0000000000000000",
50789 => "0000000000000000",50790 => "0000000000000000",
50791 => "0000000000000000",50792 => "0000000000000000",
50793 => "0000000000000000",50794 => "0000000000000000",
50795 => "0000000000000000",50796 => "0000000000000000",
50797 => "0000000000000000",50798 => "0000000000000000",
50799 => "0000000000000000",50800 => "0000000000000000",
50801 => "0000000000000000",50802 => "0000000000000000",
50803 => "0000000000000000",50804 => "0000000000000000",
50805 => "0000000000000000",50806 => "0000000000000000",
50807 => "0000000000000000",50808 => "0000000000000000",
50809 => "0000000000000000",50810 => "0000000000000000",
50811 => "0000000000000000",50812 => "0000000000000000",
50813 => "0000000000000000",50814 => "0000000000000000",
50815 => "0000000000000000",50816 => "0000000000000000",
50817 => "0000000000000000",50818 => "0000000000000000",
50819 => "0000000000000000",50820 => "0000000000000000",
50821 => "0000000000000000",50822 => "0000000000000000",
50823 => "0000000000000000",50824 => "0000000000000000",
50825 => "0000000000000000",50826 => "0000000000000000",
50827 => "0000000000000000",50828 => "0000000000000000",
50829 => "0000000000000000",50830 => "0000000000000000",
50831 => "0000000000000000",50832 => "0000000000000000",
50833 => "0000000000000000",50834 => "0000000000000000",
50835 => "0000000000000000",50836 => "0000000000000000",
50837 => "0000000000000000",50838 => "0000000000000000",
50839 => "0000000000000000",50840 => "0000000000000000",
50841 => "0000000000000000",50842 => "0000000000000000",
50843 => "0000000000000000",50844 => "0000000000000000",
50845 => "0000000000000000",50846 => "0000000000000000",
50847 => "0000000000000000",50848 => "0000000000000000",
50849 => "0000000000000000",50850 => "0000000000000000",
50851 => "0000000000000000",50852 => "0000000000000000",
50853 => "0000000000000000",50854 => "0000000000000000",
50855 => "0000000000000000",50856 => "0000000000000000",
50857 => "0000000000000000",50858 => "0000000000000000",
50859 => "0000000000000000",50860 => "0000000000000000",
50861 => "0000000000000000",50862 => "0000000000000000",
50863 => "0000000000000000",50864 => "0000000000000000",
50865 => "0000000000000000",50866 => "0000000000000000",
50867 => "0000000000000000",50868 => "0000000000000000",
50869 => "0000000000000000",50870 => "0000000000000000",
50871 => "0000000000000000",50872 => "0000000000000000",
50873 => "0000000000000000",50874 => "0000000000000000",
50875 => "0000000000000000",50876 => "0000000000000000",
50877 => "0000000000000000",50878 => "0000000000000000",
50879 => "0000000000000000",50880 => "0000000000000000",
50881 => "0000000000000000",50882 => "0000000000000000",
50883 => "0000000000000000",50884 => "0000000000000000",
50885 => "0000000000000000",50886 => "0000000000000000",
50887 => "0000000000000000",50888 => "0000000000000000",
50889 => "0000000000000000",50890 => "0000000000000000",
50891 => "0000000000000000",50892 => "0000000000000000",
50893 => "0000000000000000",50894 => "0000000000000000",
50895 => "0000000000000000",50896 => "0000000000000000",
50897 => "0000000000000000",50898 => "0000000000000000",
50899 => "0000000000000000",50900 => "0000000000000000",
50901 => "0000000000000000",50902 => "0000000000000000",
50903 => "0000000000000000",50904 => "0000000000000000",
50905 => "0000000000000000",50906 => "0000000000000000",
50907 => "0000000000000000",50908 => "0000000000000000",
50909 => "0000000000000000",50910 => "0000000000000000",
50911 => "0000000000000000",50912 => "0000000000000000",
50913 => "0000000000000000",50914 => "0000000000000000",
50915 => "0000000000000000",50916 => "0000000000000000",
50917 => "0000000000000000",50918 => "0000000000000000",
50919 => "0000000000000000",50920 => "0000000000000000",
50921 => "0000000000000000",50922 => "0000000000000000",
50923 => "0000000000000000",50924 => "0000000000000000",
50925 => "0000000000000000",50926 => "0000000000000000",
50927 => "0000000000000000",50928 => "0000000000000000",
50929 => "0000000000000000",50930 => "0000000000000000",
50931 => "0000000000000000",50932 => "0000000000000000",
50933 => "0000000000000000",50934 => "0000000000000000",
50935 => "0000000000000000",50936 => "0000000000000000",
50937 => "0000000000000000",50938 => "0000000000000000",
50939 => "0000000000000000",50940 => "0000000000000000",
50941 => "0000000000000000",50942 => "0000000000000000",
50943 => "0000000000000000",50944 => "0000000000000000",
50945 => "0000000000000000",50946 => "0000000000000000",
50947 => "0000000000000000",50948 => "0000000000000000",
50949 => "0000000000000000",50950 => "0000000000000000",
50951 => "0000000000000000",50952 => "0000000000000000",
50953 => "0000000000000000",50954 => "0000000000000000",
50955 => "0000000000000000",50956 => "0000000000000000",
50957 => "0000000000000000",50958 => "0000000000000000",
50959 => "0000000000000000",50960 => "0000000000000000",
50961 => "0000000000000000",50962 => "0000000000000000",
50963 => "0000000000000000",50964 => "0000000000000000",
50965 => "0000000000000000",50966 => "0000000000000000",
50967 => "0000000000000000",50968 => "0000000000000000",
50969 => "0000000000000000",50970 => "0000000000000000",
50971 => "0000000000000000",50972 => "0000000000000000",
50973 => "0000000000000000",50974 => "0000000000000000",
50975 => "0000000000000000",50976 => "0000000000000000",
50977 => "0000000000000000",50978 => "0000000000000000",
50979 => "0000000000000000",50980 => "0000000000000000",
50981 => "0000000000000000",50982 => "0000000000000000",
50983 => "0000000000000000",50984 => "0000000000000000",
50985 => "0000000000000000",50986 => "0000000000000000",
50987 => "0000000000000000",50988 => "0000000000000000",
50989 => "0000000000000000",50990 => "0000000000000000",
50991 => "0000000000000000",50992 => "0000000000000000",
50993 => "0000000000000000",50994 => "0000000000000000",
50995 => "0000000000000000",50996 => "0000000000000000",
50997 => "0000000000000000",50998 => "0000000000000000",
50999 => "0000000000000000",51000 => "0000000000000000",
51001 => "0000000000000000",51002 => "0000000000000000",
51003 => "0000000000000000",51004 => "0000000000000000",
51005 => "0000000000000000",51006 => "0000000000000000",
51007 => "0000000000000000",51008 => "0000000000000000",
51009 => "0000000000000000",51010 => "0000000000000000",
51011 => "0000000000000000",51012 => "0000000000000000",
51013 => "0000000000000000",51014 => "0000000000000000",
51015 => "0000000000000000",51016 => "0000000000000000",
51017 => "0000000000000000",51018 => "0000000000000000",
51019 => "0000000000000000",51020 => "0000000000000000",
51021 => "0000000000000000",51022 => "0000000000000000",
51023 => "0000000000000000",51024 => "0000000000000000",
51025 => "0000000000000000",51026 => "0000000000000000",
51027 => "0000000000000000",51028 => "0000000000000000",
51029 => "0000000000000000",51030 => "0000000000000000",
51031 => "0000000000000000",51032 => "0000000000000000",
51033 => "0000000000000000",51034 => "0000000000000000",
51035 => "0000000000000000",51036 => "0000000000000000",
51037 => "0000000000000000",51038 => "0000000000000000",
51039 => "0000000000000000",51040 => "0000000000000000",
51041 => "0000000000000000",51042 => "0000000000000000",
51043 => "0000000000000000",51044 => "0000000000000000",
51045 => "0000000000000000",51046 => "0000000000000000",
51047 => "0000000000000000",51048 => "0000000000000000",
51049 => "0000000000000000",51050 => "0000000000000000",
51051 => "0000000000000000",51052 => "0000000000000000",
51053 => "0000000000000000",51054 => "0000000000000000",
51055 => "0000000000000000",51056 => "0000000000000000",
51057 => "0000000000000000",51058 => "0000000000000000",
51059 => "0000000000000000",51060 => "0000000000000000",
51061 => "0000000000000000",51062 => "0000000000000000",
51063 => "0000000000000000",51064 => "0000000000000000",
51065 => "0000000000000000",51066 => "0000000000000000",
51067 => "0000000000000000",51068 => "0000000000000000",
51069 => "0000000000000000",51070 => "0000000000000000",
51071 => "0000000000000000",51072 => "0000000000000000",
51073 => "0000000000000000",51074 => "0000000000000000",
51075 => "0000000000000000",51076 => "0000000000000000",
51077 => "0000000000000000",51078 => "0000000000000000",
51079 => "0000000000000000",51080 => "0000000000000000",
51081 => "0000000000000000",51082 => "0000000000000000",
51083 => "0000000000000000",51084 => "0000000000000000",
51085 => "0000000000000000",51086 => "0000000000000000",
51087 => "0000000000000000",51088 => "0000000000000000",
51089 => "0000000000000000",51090 => "0000000000000000",
51091 => "0000000000000000",51092 => "0000000000000000",
51093 => "0000000000000000",51094 => "0000000000000000",
51095 => "0000000000000000",51096 => "0000000000000000",
51097 => "0000000000000000",51098 => "0000000000000000",
51099 => "0000000000000000",51100 => "0000000000000000",
51101 => "0000000000000000",51102 => "0000000000000000",
51103 => "0000000000000000",51104 => "0000000000000000",
51105 => "0000000000000000",51106 => "0000000000000000",
51107 => "0000000000000000",51108 => "0000000000000000",
51109 => "0000000000000000",51110 => "0000000000000000",
51111 => "0000000000000000",51112 => "0000000000000000",
51113 => "0000000000000000",51114 => "0000000000000000",
51115 => "0000000000000000",51116 => "0000000000000000",
51117 => "0000000000000000",51118 => "0000000000000000",
51119 => "0000000000000000",51120 => "0000000000000000",
51121 => "0000000000000000",51122 => "0000000000000000",
51123 => "0000000000000000",51124 => "0000000000000000",
51125 => "0000000000000000",51126 => "0000000000000000",
51127 => "0000000000000000",51128 => "0000000000000000",
51129 => "0000000000000000",51130 => "0000000000000000",
51131 => "0000000000000000",51132 => "0000000000000000",
51133 => "0000000000000000",51134 => "0000000000000000",
51135 => "0000000000000000",51136 => "0000000000000000",
51137 => "0000000000000000",51138 => "0000000000000000",
51139 => "0000000000000000",51140 => "0000000000000000",
51141 => "0000000000000000",51142 => "0000000000000000",
51143 => "0000000000000000",51144 => "0000000000000000",
51145 => "0000000000000000",51146 => "0000000000000000",
51147 => "0000000000000000",51148 => "0000000000000000",
51149 => "0000000000000000",51150 => "0000000000000000",
51151 => "0000000000000000",51152 => "0000000000000000",
51153 => "0000000000000000",51154 => "0000000000000000",
51155 => "0000000000000000",51156 => "0000000000000000",
51157 => "0000000000000000",51158 => "0000000000000000",
51159 => "0000000000000000",51160 => "0000000000000000",
51161 => "0000000000000000",51162 => "0000000000000000",
51163 => "0000000000000000",51164 => "0000000000000000",
51165 => "0000000000000000",51166 => "0000000000000000",
51167 => "0000000000000000",51168 => "0000000000000000",
51169 => "0000000000000000",51170 => "0000000000000000",
51171 => "0000000000000000",51172 => "0000000000000000",
51173 => "0000000000000000",51174 => "0000000000000000",
51175 => "0000000000000000",51176 => "0000000000000000",
51177 => "0000000000000000",51178 => "0000000000000000",
51179 => "0000000000000000",51180 => "0000000000000000",
51181 => "0000000000000000",51182 => "0000000000000000",
51183 => "0000000000000000",51184 => "0000000000000000",
51185 => "0000000000000000",51186 => "0000000000000000",
51187 => "0000000000000000",51188 => "0000000000000000",
51189 => "0000000000000000",51190 => "0000000000000000",
51191 => "0000000000000000",51192 => "0000000000000000",
51193 => "0000000000000000",51194 => "0000000000000000",
51195 => "0000000000000000",51196 => "0000000000000000",
51197 => "0000000000000000",51198 => "0000000000000000",
51199 => "0000000000000000",51200 => "0000000000000000",
51201 => "0000000000000000",51202 => "0000000000000000",
51203 => "0000000000000000",51204 => "0000000000000000",
51205 => "0000000000000000",51206 => "0000000000000000",
51207 => "0000000000000000",51208 => "0000000000000000",
51209 => "0000000000000000",51210 => "0000000000000000",
51211 => "0000000000000000",51212 => "0000000000000000",
51213 => "0000000000000000",51214 => "0000000000000000",
51215 => "0000000000000000",51216 => "0000000000000000",
51217 => "0000000000000000",51218 => "0000000000000000",
51219 => "0000000000000000",51220 => "0000000000000000",
51221 => "0000000000000000",51222 => "0000000000000000",
51223 => "0000000000000000",51224 => "0000000000000000",
51225 => "0000000000000000",51226 => "0000000000000000",
51227 => "0000000000000000",51228 => "0000000000000000",
51229 => "0000000000000000",51230 => "0000000000000000",
51231 => "0000000000000000",51232 => "0000000000000000",
51233 => "0000000000000000",51234 => "0000000000000000",
51235 => "0000000000000000",51236 => "0000000000000000",
51237 => "0000000000000000",51238 => "0000000000000000",
51239 => "0000000000000000",51240 => "0000000000000000",
51241 => "0000000000000000",51242 => "0000000000000000",
51243 => "0000000000000000",51244 => "0000000000000000",
51245 => "0000000000000000",51246 => "0000000000000000",
51247 => "0000000000000000",51248 => "0000000000000000",
51249 => "0000000000000000",51250 => "0000000000000000",
51251 => "0000000000000000",51252 => "0000000000000000",
51253 => "0000000000000000",51254 => "0000000000000000",
51255 => "0000000000000000",51256 => "0000000000000000",
51257 => "0000000000000000",51258 => "0000000000000000",
51259 => "0000000000000000",51260 => "0000000000000000",
51261 => "0000000000000000",51262 => "0000000000000000",
51263 => "0000000000000000",51264 => "0000000000000000",
51265 => "0000000000000000",51266 => "0000000000000000",
51267 => "0000000000000000",51268 => "0000000000000000",
51269 => "0000000000000000",51270 => "0000000000000000",
51271 => "0000000000000000",51272 => "0000000000000000",
51273 => "0000000000000000",51274 => "0000000000000000",
51275 => "0000000000000000",51276 => "0000000000000000",
51277 => "0000000000000000",51278 => "0000000000000000",
51279 => "0000000000000000",51280 => "0000000000000000",
51281 => "0000000000000000",51282 => "0000000000000000",
51283 => "0000000000000000",51284 => "0000000000000000",
51285 => "0000000000000000",51286 => "0000000000000000",
51287 => "0000000000000000",51288 => "0000000000000000",
51289 => "0000000000000000",51290 => "0000000000000000",
51291 => "0000000000000000",51292 => "0000000000000000",
51293 => "0000000000000000",51294 => "0000000000000000",
51295 => "0000000000000000",51296 => "0000000000000000",
51297 => "0000000000000000",51298 => "0000000000000000",
51299 => "0000000000000000",51300 => "0000000000000000",
51301 => "0000000000000000",51302 => "0000000000000000",
51303 => "0000000000000000",51304 => "0000000000000000",
51305 => "0000000000000000",51306 => "0000000000000000",
51307 => "0000000000000000",51308 => "0000000000000000",
51309 => "0000000000000000",51310 => "0000000000000000",
51311 => "0000000000000000",51312 => "0000000000000000",
51313 => "0000000000000000",51314 => "0000000000000000",
51315 => "0000000000000000",51316 => "0000000000000000",
51317 => "0000000000000000",51318 => "0000000000000000",
51319 => "0000000000000000",51320 => "0000000000000000",
51321 => "0000000000000000",51322 => "0000000000000000",
51323 => "0000000000000000",51324 => "0000000000000000",
51325 => "0000000000000000",51326 => "0000000000000000",
51327 => "0000000000000000",51328 => "0000000000000000",
51329 => "0000000000000000",51330 => "0000000000000000",
51331 => "0000000000000000",51332 => "0000000000000000",
51333 => "0000000000000000",51334 => "0000000000000000",
51335 => "0000000000000000",51336 => "0000000000000000",
51337 => "0000000000000000",51338 => "0000000000000000",
51339 => "0000000000000000",51340 => "0000000000000000",
51341 => "0000000000000000",51342 => "0000000000000000",
51343 => "0000000000000000",51344 => "0000000000000000",
51345 => "0000000000000000",51346 => "0000000000000000",
51347 => "0000000000000000",51348 => "0000000000000000",
51349 => "0000000000000000",51350 => "0000000000000000",
51351 => "0000000000000000",51352 => "0000000000000000",
51353 => "0000000000000000",51354 => "0000000000000000",
51355 => "0000000000000000",51356 => "0000000000000000",
51357 => "0000000000000000",51358 => "0000000000000000",
51359 => "0000000000000000",51360 => "0000000000000000",
51361 => "0000000000000000",51362 => "0000000000000000",
51363 => "0000000000000000",51364 => "0000000000000000",
51365 => "0000000000000000",51366 => "0000000000000000",
51367 => "0000000000000000",51368 => "0000000000000000",
51369 => "0000000000000000",51370 => "0000000000000000",
51371 => "0000000000000000",51372 => "0000000000000000",
51373 => "0000000000000000",51374 => "0000000000000000",
51375 => "0000000000000000",51376 => "0000000000000000",
51377 => "0000000000000000",51378 => "0000000000000000",
51379 => "0000000000000000",51380 => "0000000000000000",
51381 => "0000000000000000",51382 => "0000000000000000",
51383 => "0000000000000000",51384 => "0000000000000000",
51385 => "0000000000000000",51386 => "0000000000000000",
51387 => "0000000000000000",51388 => "0000000000000000",
51389 => "0000000000000000",51390 => "0000000000000000",
51391 => "0000000000000000",51392 => "0000000000000000",
51393 => "0000000000000000",51394 => "0000000000000000",
51395 => "0000000000000000",51396 => "0000000000000000",
51397 => "0000000000000000",51398 => "0000000000000000",
51399 => "0000000000000000",51400 => "0000000000000000",
51401 => "0000000000000000",51402 => "0000000000000000",
51403 => "0000000000000000",51404 => "0000000000000000",
51405 => "0000000000000000",51406 => "0000000000000000",
51407 => "0000000000000000",51408 => "0000000000000000",
51409 => "0000000000000000",51410 => "0000000000000000",
51411 => "0000000000000000",51412 => "0000000000000000",
51413 => "0000000000000000",51414 => "0000000000000000",
51415 => "0000000000000000",51416 => "0000000000000000",
51417 => "0000000000000000",51418 => "0000000000000000",
51419 => "0000000000000000",51420 => "0000000000000000",
51421 => "0000000000000000",51422 => "0000000000000000",
51423 => "0000000000000000",51424 => "0000000000000000",
51425 => "0000000000000000",51426 => "0000000000000000",
51427 => "0000000000000000",51428 => "0000000000000000",
51429 => "0000000000000000",51430 => "0000000000000000",
51431 => "0000000000000000",51432 => "0000000000000000",
51433 => "0000000000000000",51434 => "0000000000000000",
51435 => "0000000000000000",51436 => "0000000000000000",
51437 => "0000000000000000",51438 => "0000000000000000",
51439 => "0000000000000000",51440 => "0000000000000000",
51441 => "0000000000000000",51442 => "0000000000000000",
51443 => "0000000000000000",51444 => "0000000000000000",
51445 => "0000000000000000",51446 => "0000000000000000",
51447 => "0000000000000000",51448 => "0000000000000000",
51449 => "0000000000000000",51450 => "0000000000000000",
51451 => "0000000000000000",51452 => "0000000000000000",
51453 => "0000000000000000",51454 => "0000000000000000",
51455 => "0000000000000000",51456 => "0000000000000000",
51457 => "0000000000000000",51458 => "0000000000000000",
51459 => "0000000000000000",51460 => "0000000000000000",
51461 => "0000000000000000",51462 => "0000000000000000",
51463 => "0000000000000000",51464 => "0000000000000000",
51465 => "0000000000000000",51466 => "0000000000000000",
51467 => "0000000000000000",51468 => "0000000000000000",
51469 => "0000000000000000",51470 => "0000000000000000",
51471 => "0000000000000000",51472 => "0000000000000000",
51473 => "0000000000000000",51474 => "0000000000000000",
51475 => "0000000000000000",51476 => "0000000000000000",
51477 => "0000000000000000",51478 => "0000000000000000",
51479 => "0000000000000000",51480 => "0000000000000000",
51481 => "0000000000000000",51482 => "0000000000000000",
51483 => "0000000000000000",51484 => "0000000000000000",
51485 => "0000000000000000",51486 => "0000000000000000",
51487 => "0000000000000000",51488 => "0000000000000000",
51489 => "0000000000000000",51490 => "0000000000000000",
51491 => "0000000000000000",51492 => "0000000000000000",
51493 => "0000000000000000",51494 => "0000000000000000",
51495 => "0000000000000000",51496 => "0000000000000000",
51497 => "0000000000000000",51498 => "0000000000000000",
51499 => "0000000000000000",51500 => "0000000000000000",
51501 => "0000000000000000",51502 => "0000000000000000",
51503 => "0000000000000000",51504 => "0000000000000000",
51505 => "0000000000000000",51506 => "0000000000000000",
51507 => "0000000000000000",51508 => "0000000000000000",
51509 => "0000000000000000",51510 => "0000000000000000",
51511 => "0000000000000000",51512 => "0000000000000000",
51513 => "0000000000000000",51514 => "0000000000000000",
51515 => "0000000000000000",51516 => "0000000000000000",
51517 => "0000000000000000",51518 => "0000000000000000",
51519 => "0000000000000000",51520 => "0000000000000000",
51521 => "0000000000000000",51522 => "0000000000000000",
51523 => "0000000000000000",51524 => "0000000000000000",
51525 => "0000000000000000",51526 => "0000000000000000",
51527 => "0000000000000000",51528 => "0000000000000000",
51529 => "0000000000000000",51530 => "0000000000000000",
51531 => "0000000000000000",51532 => "0000000000000000",
51533 => "0000000000000000",51534 => "0000000000000000",
51535 => "0000000000000000",51536 => "0000000000000000",
51537 => "0000000000000000",51538 => "0000000000000000",
51539 => "0000000000000000",51540 => "0000000000000000",
51541 => "0000000000000000",51542 => "0000000000000000",
51543 => "0000000000000000",51544 => "0000000000000000",
51545 => "0000000000000000",51546 => "0000000000000000",
51547 => "0000000000000000",51548 => "0000000000000000",
51549 => "0000000000000000",51550 => "0000000000000000",
51551 => "0000000000000000",51552 => "0000000000000000",
51553 => "0000000000000000",51554 => "0000000000000000",
51555 => "0000000000000000",51556 => "0000000000000000",
51557 => "0000000000000000",51558 => "0000000000000000",
51559 => "0000000000000000",51560 => "0000000000000000",
51561 => "0000000000000000",51562 => "0000000000000000",
51563 => "0000000000000000",51564 => "0000000000000000",
51565 => "0000000000000000",51566 => "0000000000000000",
51567 => "0000000000000000",51568 => "0000000000000000",
51569 => "0000000000000000",51570 => "0000000000000000",
51571 => "0000000000000000",51572 => "0000000000000000",
51573 => "0000000000000000",51574 => "0000000000000000",
51575 => "0000000000000000",51576 => "0000000000000000",
51577 => "0000000000000000",51578 => "0000000000000000",
51579 => "0000000000000000",51580 => "0000000000000000",
51581 => "0000000000000000",51582 => "0000000000000000",
51583 => "0000000000000000",51584 => "0000000000000000",
51585 => "0000000000000000",51586 => "0000000000000000",
51587 => "0000000000000000",51588 => "0000000000000000",
51589 => "0000000000000000",51590 => "0000000000000000",
51591 => "0000000000000000",51592 => "0000000000000000",
51593 => "0000000000000000",51594 => "0000000000000000",
51595 => "0000000000000000",51596 => "0000000000000000",
51597 => "0000000000000000",51598 => "0000000000000000",
51599 => "0000000000000000",51600 => "0000000000000000",
51601 => "0000000000000000",51602 => "0000000000000000",
51603 => "0000000000000000",51604 => "0000000000000000",
51605 => "0000000000000000",51606 => "0000000000000000",
51607 => "0000000000000000",51608 => "0000000000000000",
51609 => "0000000000000000",51610 => "0000000000000000",
51611 => "0000000000000000",51612 => "0000000000000000",
51613 => "0000000000000000",51614 => "0000000000000000",
51615 => "0000000000000000",51616 => "0000000000000000",
51617 => "0000000000000000",51618 => "0000000000000000",
51619 => "0000000000000000",51620 => "0000000000000000",
51621 => "0000000000000000",51622 => "0000000000000000",
51623 => "0000000000000000",51624 => "0000000000000000",
51625 => "0000000000000000",51626 => "0000000000000000",
51627 => "0000000000000000",51628 => "0000000000000000",
51629 => "0000000000000000",51630 => "0000000000000000",
51631 => "0000000000000000",51632 => "0000000000000000",
51633 => "0000000000000000",51634 => "0000000000000000",
51635 => "0000000000000000",51636 => "0000000000000000",
51637 => "0000000000000000",51638 => "0000000000000000",
51639 => "0000000000000000",51640 => "0000000000000000",
51641 => "0000000000000000",51642 => "0000000000000000",
51643 => "0000000000000000",51644 => "0000000000000000",
51645 => "0000000000000000",51646 => "0000000000000000",
51647 => "0000000000000000",51648 => "0000000000000000",
51649 => "0000000000000000",51650 => "0000000000000000",
51651 => "0000000000000000",51652 => "0000000000000000",
51653 => "0000000000000000",51654 => "0000000000000000",
51655 => "0000000000000000",51656 => "0000000000000000",
51657 => "0000000000000000",51658 => "0000000000000000",
51659 => "0000000000000000",51660 => "0000000000000000",
51661 => "0000000000000000",51662 => "0000000000000000",
51663 => "0000000000000000",51664 => "0000000000000000",
51665 => "0000000000000000",51666 => "0000000000000000",
51667 => "0000000000000000",51668 => "0000000000000000",
51669 => "0000000000000000",51670 => "0000000000000000",
51671 => "0000000000000000",51672 => "0000000000000000",
51673 => "0000000000000000",51674 => "0000000000000000",
51675 => "0000000000000000",51676 => "0000000000000000",
51677 => "0000000000000000",51678 => "0000000000000000",
51679 => "0000000000000000",51680 => "0000000000000000",
51681 => "0000000000000000",51682 => "0000000000000000",
51683 => "0000000000000000",51684 => "0000000000000000",
51685 => "0000000000000000",51686 => "0000000000000000",
51687 => "0000000000000000",51688 => "0000000000000000",
51689 => "0000000000000000",51690 => "0000000000000000",
51691 => "0000000000000000",51692 => "0000000000000000",
51693 => "0000000000000000",51694 => "0000000000000000",
51695 => "0000000000000000",51696 => "0000000000000000",
51697 => "0000000000000000",51698 => "0000000000000000",
51699 => "0000000000000000",51700 => "0000000000000000",
51701 => "0000000000000000",51702 => "0000000000000000",
51703 => "0000000000000000",51704 => "0000000000000000",
51705 => "0000000000000000",51706 => "0000000000000000",
51707 => "0000000000000000",51708 => "0000000000000000",
51709 => "0000000000000000",51710 => "0000000000000000",
51711 => "0000000000000000",51712 => "0000000000000000",
51713 => "0000000000000000",51714 => "0000000000000000",
51715 => "0000000000000000",51716 => "0000000000000000",
51717 => "0000000000000000",51718 => "0000000000000000",
51719 => "0000000000000000",51720 => "0000000000000000",
51721 => "0000000000000000",51722 => "0000000000000000",
51723 => "0000000000000000",51724 => "0000000000000000",
51725 => "0000000000000000",51726 => "0000000000000000",
51727 => "0000000000000000",51728 => "0000000000000000",
51729 => "0000000000000000",51730 => "0000000000000000",
51731 => "0000000000000000",51732 => "0000000000000000",
51733 => "0000000000000000",51734 => "0000000000000000",
51735 => "0000000000000000",51736 => "0000000000000000",
51737 => "0000000000000000",51738 => "0000000000000000",
51739 => "0000000000000000",51740 => "0000000000000000",
51741 => "0000000000000000",51742 => "0000000000000000",
51743 => "0000000000000000",51744 => "0000000000000000",
51745 => "0000000000000000",51746 => "0000000000000000",
51747 => "0000000000000000",51748 => "0000000000000000",
51749 => "0000000000000000",51750 => "0000000000000000",
51751 => "0000000000000000",51752 => "0000000000000000",
51753 => "0000000000000000",51754 => "0000000000000000",
51755 => "0000000000000000",51756 => "0000000000000000",
51757 => "0000000000000000",51758 => "0000000000000000",
51759 => "0000000000000000",51760 => "0000000000000000",
51761 => "0000000000000000",51762 => "0000000000000000",
51763 => "0000000000000000",51764 => "0000000000000000",
51765 => "0000000000000000",51766 => "0000000000000000",
51767 => "0000000000000000",51768 => "0000000000000000",
51769 => "0000000000000000",51770 => "0000000000000000",
51771 => "0000000000000000",51772 => "0000000000000000",
51773 => "0000000000000000",51774 => "0000000000000000",
51775 => "0000000000000000",51776 => "0000000000000000",
51777 => "0000000000000000",51778 => "0000000000000000",
51779 => "0000000000000000",51780 => "0000000000000000",
51781 => "0000000000000000",51782 => "0000000000000000",
51783 => "0000000000000000",51784 => "0000000000000000",
51785 => "0000000000000000",51786 => "0000000000000000",
51787 => "0000000000000000",51788 => "0000000000000000",
51789 => "0000000000000000",51790 => "0000000000000000",
51791 => "0000000000000000",51792 => "0000000000000000",
51793 => "0000000000000000",51794 => "0000000000000000",
51795 => "0000000000000000",51796 => "0000000000000000",
51797 => "0000000000000000",51798 => "0000000000000000",
51799 => "0000000000000000",51800 => "0000000000000000",
51801 => "0000000000000000",51802 => "0000000000000000",
51803 => "0000000000000000",51804 => "0000000000000000",
51805 => "0000000000000000",51806 => "0000000000000000",
51807 => "0000000000000000",51808 => "0000000000000000",
51809 => "0000000000000000",51810 => "0000000000000000",
51811 => "0000000000000000",51812 => "0000000000000000",
51813 => "0000000000000000",51814 => "0000000000000000",
51815 => "0000000000000000",51816 => "0000000000000000",
51817 => "0000000000000000",51818 => "0000000000000000",
51819 => "0000000000000000",51820 => "0000000000000000",
51821 => "0000000000000000",51822 => "0000000000000000",
51823 => "0000000000000000",51824 => "0000000000000000",
51825 => "0000000000000000",51826 => "0000000000000000",
51827 => "0000000000000000",51828 => "0000000000000000",
51829 => "0000000000000000",51830 => "0000000000000000",
51831 => "0000000000000000",51832 => "0000000000000000",
51833 => "0000000000000000",51834 => "0000000000000000",
51835 => "0000000000000000",51836 => "0000000000000000",
51837 => "0000000000000000",51838 => "0000000000000000",
51839 => "0000000000000000",51840 => "0000000000000000",
51841 => "0000000000000000",51842 => "0000000000000000",
51843 => "0000000000000000",51844 => "0000000000000000",
51845 => "0000000000000000",51846 => "0000000000000000",
51847 => "0000000000000000",51848 => "0000000000000000",
51849 => "0000000000000000",51850 => "0000000000000000",
51851 => "0000000000000000",51852 => "0000000000000000",
51853 => "0000000000000000",51854 => "0000000000000000",
51855 => "0000000000000000",51856 => "0000000000000000",
51857 => "0000000000000000",51858 => "0000000000000000",
51859 => "0000000000000000",51860 => "0000000000000000",
51861 => "0000000000000000",51862 => "0000000000000000",
51863 => "0000000000000000",51864 => "0000000000000000",
51865 => "0000000000000000",51866 => "0000000000000000",
51867 => "0000000000000000",51868 => "0000000000000000",
51869 => "0000000000000000",51870 => "0000000000000000",
51871 => "0000000000000000",51872 => "0000000000000000",
51873 => "0000000000000000",51874 => "0000000000000000",
51875 => "0000000000000000",51876 => "0000000000000000",
51877 => "0000000000000000",51878 => "0000000000000000",
51879 => "0000000000000000",51880 => "0000000000000000",
51881 => "0000000000000000",51882 => "0000000000000000",
51883 => "0000000000000000",51884 => "0000000000000000",
51885 => "0000000000000000",51886 => "0000000000000000",
51887 => "0000000000000000",51888 => "0000000000000000",
51889 => "0000000000000000",51890 => "0000000000000000",
51891 => "0000000000000000",51892 => "0000000000000000",
51893 => "0000000000000000",51894 => "0000000000000000",
51895 => "0000000000000000",51896 => "0000000000000000",
51897 => "0000000000000000",51898 => "0000000000000000",
51899 => "0000000000000000",51900 => "0000000000000000",
51901 => "0000000000000000",51902 => "0000000000000000",
51903 => "0000000000000000",51904 => "0000000000000000",
51905 => "0000000000000000",51906 => "0000000000000000",
51907 => "0000000000000000",51908 => "0000000000000000",
51909 => "0000000000000000",51910 => "0000000000000000",
51911 => "0000000000000000",51912 => "0000000000000000",
51913 => "0000000000000000",51914 => "0000000000000000",
51915 => "0000000000000000",51916 => "0000000000000000",
51917 => "0000000000000000",51918 => "0000000000000000",
51919 => "0000000000000000",51920 => "0000000000000000",
51921 => "0000000000000000",51922 => "0000000000000000",
51923 => "0000000000000000",51924 => "0000000000000000",
51925 => "0000000000000000",51926 => "0000000000000000",
51927 => "0000000000000000",51928 => "0000000000000000",
51929 => "0000000000000000",51930 => "0000000000000000",
51931 => "0000000000000000",51932 => "0000000000000000",
51933 => "0000000000000000",51934 => "0000000000000000",
51935 => "0000000000000000",51936 => "0000000000000000",
51937 => "0000000000000000",51938 => "0000000000000000",
51939 => "0000000000000000",51940 => "0000000000000000",
51941 => "0000000000000000",51942 => "0000000000000000",
51943 => "0000000000000000",51944 => "0000000000000000",
51945 => "0000000000000000",51946 => "0000000000000000",
51947 => "0000000000000000",51948 => "0000000000000000",
51949 => "0000000000000000",51950 => "0000000000000000",
51951 => "0000000000000000",51952 => "0000000000000000",
51953 => "0000000000000000",51954 => "0000000000000000",
51955 => "0000000000000000",51956 => "0000000000000000",
51957 => "0000000000000000",51958 => "0000000000000000",
51959 => "0000000000000000",51960 => "0000000000000000",
51961 => "0000000000000000",51962 => "0000000000000000",
51963 => "0000000000000000",51964 => "0000000000000000",
51965 => "0000000000000000",51966 => "0000000000000000",
51967 => "0000000000000000",51968 => "0000000000000000",
51969 => "0000000000000000",51970 => "0000000000000000",
51971 => "0000000000000000",51972 => "0000000000000000",
51973 => "0000000000000000",51974 => "0000000000000000",
51975 => "0000000000000000",51976 => "0000000000000000",
51977 => "0000000000000000",51978 => "0000000000000000",
51979 => "0000000000000000",51980 => "0000000000000000",
51981 => "0000000000000000",51982 => "0000000000000000",
51983 => "0000000000000000",51984 => "0000000000000000",
51985 => "0000000000000000",51986 => "0000000000000000",
51987 => "0000000000000000",51988 => "0000000000000000",
51989 => "0000000000000000",51990 => "0000000000000000",
51991 => "0000000000000000",51992 => "0000000000000000",
51993 => "0000000000000000",51994 => "0000000000000000",
51995 => "0000000000000000",51996 => "0000000000000000",
51997 => "0000000000000000",51998 => "0000000000000000",
51999 => "0000000000000000",52000 => "0000000000000000",
52001 => "0000000000000000",52002 => "0000000000000000",
52003 => "0000000000000000",52004 => "0000000000000000",
52005 => "0000000000000000",52006 => "0000000000000000",
52007 => "0000000000000000",52008 => "0000000000000000",
52009 => "0000000000000000",52010 => "0000000000000000",
52011 => "0000000000000000",52012 => "0000000000000000",
52013 => "0000000000000000",52014 => "0000000000000000",
52015 => "0000000000000000",52016 => "0000000000000000",
52017 => "0000000000000000",52018 => "0000000000000000",
52019 => "0000000000000000",52020 => "0000000000000000",
52021 => "0000000000000000",52022 => "0000000000000000",
52023 => "0000000000000000",52024 => "0000000000000000",
52025 => "0000000000000000",52026 => "0000000000000000",
52027 => "0000000000000000",52028 => "0000000000000000",
52029 => "0000000000000000",52030 => "0000000000000000",
52031 => "0000000000000000",52032 => "0000000000000000",
52033 => "0000000000000000",52034 => "0000000000000000",
52035 => "0000000000000000",52036 => "0000000000000000",
52037 => "0000000000000000",52038 => "0000000000000000",
52039 => "0000000000000000",52040 => "0000000000000000",
52041 => "0000000000000000",52042 => "0000000000000000",
52043 => "0000000000000000",52044 => "0000000000000000",
52045 => "0000000000000000",52046 => "0000000000000000",
52047 => "0000000000000000",52048 => "0000000000000000",
52049 => "0000000000000000",52050 => "0000000000000000",
52051 => "0000000000000000",52052 => "0000000000000000",
52053 => "0000000000000000",52054 => "0000000000000000",
52055 => "0000000000000000",52056 => "0000000000000000",
52057 => "0000000000000000",52058 => "0000000000000000",
52059 => "0000000000000000",52060 => "0000000000000000",
52061 => "0000000000000000",52062 => "0000000000000000",
52063 => "0000000000000000",52064 => "0000000000000000",
52065 => "0000000000000000",52066 => "0000000000000000",
52067 => "0000000000000000",52068 => "0000000000000000",
52069 => "0000000000000000",52070 => "0000000000000000",
52071 => "0000000000000000",52072 => "0000000000000000",
52073 => "0000000000000000",52074 => "0000000000000000",
52075 => "0000000000000000",52076 => "0000000000000000",
52077 => "0000000000000000",52078 => "0000000000000000",
52079 => "0000000000000000",52080 => "0000000000000000",
52081 => "0000000000000000",52082 => "0000000000000000",
52083 => "0000000000000000",52084 => "0000000000000000",
52085 => "0000000000000000",52086 => "0000000000000000",
52087 => "0000000000000000",52088 => "0000000000000000",
52089 => "0000000000000000",52090 => "0000000000000000",
52091 => "0000000000000000",52092 => "0000000000000000",
52093 => "0000000000000000",52094 => "0000000000000000",
52095 => "0000000000000000",52096 => "0000000000000000",
52097 => "0000000000000000",52098 => "0000000000000000",
52099 => "0000000000000000",52100 => "0000000000000000",
52101 => "0000000000000000",52102 => "0000000000000000",
52103 => "0000000000000000",52104 => "0000000000000000",
52105 => "0000000000000000",52106 => "0000000000000000",
52107 => "0000000000000000",52108 => "0000000000000000",
52109 => "0000000000000000",52110 => "0000000000000000",
52111 => "0000000000000000",52112 => "0000000000000000",
52113 => "0000000000000000",52114 => "0000000000000000",
52115 => "0000000000000000",52116 => "0000000000000000",
52117 => "0000000000000000",52118 => "0000000000000000",
52119 => "0000000000000000",52120 => "0000000000000000",
52121 => "0000000000000000",52122 => "0000000000000000",
52123 => "0000000000000000",52124 => "0000000000000000",
52125 => "0000000000000000",52126 => "0000000000000000",
52127 => "0000000000000000",52128 => "0000000000000000",
52129 => "0000000000000000",52130 => "0000000000000000",
52131 => "0000000000000000",52132 => "0000000000000000",
52133 => "0000000000000000",52134 => "0000000000000000",
52135 => "0000000000000000",52136 => "0000000000000000",
52137 => "0000000000000000",52138 => "0000000000000000",
52139 => "0000000000000000",52140 => "0000000000000000",
52141 => "0000000000000000",52142 => "0000000000000000",
52143 => "0000000000000000",52144 => "0000000000000000",
52145 => "0000000000000000",52146 => "0000000000000000",
52147 => "0000000000000000",52148 => "0000000000000000",
52149 => "0000000000000000",52150 => "0000000000000000",
52151 => "0000000000000000",52152 => "0000000000000000",
52153 => "0000000000000000",52154 => "0000000000000000",
52155 => "0000000000000000",52156 => "0000000000000000",
52157 => "0000000000000000",52158 => "0000000000000000",
52159 => "0000000000000000",52160 => "0000000000000000",
52161 => "0000000000000000",52162 => "0000000000000000",
52163 => "0000000000000000",52164 => "0000000000000000",
52165 => "0000000000000000",52166 => "0000000000000000",
52167 => "0000000000000000",52168 => "0000000000000000",
52169 => "0000000000000000",52170 => "0000000000000000",
52171 => "0000000000000000",52172 => "0000000000000000",
52173 => "0000000000000000",52174 => "0000000000000000",
52175 => "0000000000000000",52176 => "0000000000000000",
52177 => "0000000000000000",52178 => "0000000000000000",
52179 => "0000000000000000",52180 => "0000000000000000",
52181 => "0000000000000000",52182 => "0000000000000000",
52183 => "0000000000000000",52184 => "0000000000000000",
52185 => "0000000000000000",52186 => "0000000000000000",
52187 => "0000000000000000",52188 => "0000000000000000",
52189 => "0000000000000000",52190 => "0000000000000000",
52191 => "0000000000000000",52192 => "0000000000000000",
52193 => "0000000000000000",52194 => "0000000000000000",
52195 => "0000000000000000",52196 => "0000000000000000",
52197 => "0000000000000000",52198 => "0000000000000000",
52199 => "0000000000000000",52200 => "0000000000000000",
52201 => "0000000000000000",52202 => "0000000000000000",
52203 => "0000000000000000",52204 => "0000000000000000",
52205 => "0000000000000000",52206 => "0000000000000000",
52207 => "0000000000000000",52208 => "0000000000000000",
52209 => "0000000000000000",52210 => "0000000000000000",
52211 => "0000000000000000",52212 => "0000000000000000",
52213 => "0000000000000000",52214 => "0000000000000000",
52215 => "0000000000000000",52216 => "0000000000000000",
52217 => "0000000000000000",52218 => "0000000000000000",
52219 => "0000000000000000",52220 => "0000000000000000",
52221 => "0000000000000000",52222 => "0000000000000000",
52223 => "0000000000000000",52224 => "0000000000000000",
52225 => "0000000000000000",52226 => "0000000000000000",
52227 => "0000000000000000",52228 => "0000000000000000",
52229 => "0000000000000000",52230 => "0000000000000000",
52231 => "0000000000000000",52232 => "0000000000000000",
52233 => "0000000000000000",52234 => "0000000000000000",
52235 => "0000000000000000",52236 => "0000000000000000",
52237 => "0000000000000000",52238 => "0000000000000000",
52239 => "0000000000000000",52240 => "0000000000000000",
52241 => "0000000000000000",52242 => "0000000000000000",
52243 => "0000000000000000",52244 => "0000000000000000",
52245 => "0000000000000000",52246 => "0000000000000000",
52247 => "0000000000000000",52248 => "0000000000000000",
52249 => "0000000000000000",52250 => "0000000000000000",
52251 => "0000000000000000",52252 => "0000000000000000",
52253 => "0000000000000000",52254 => "0000000000000000",
52255 => "0000000000000000",52256 => "0000000000000000",
52257 => "0000000000000000",52258 => "0000000000000000",
52259 => "0000000000000000",52260 => "0000000000000000",
52261 => "0000000000000000",52262 => "0000000000000000",
52263 => "0000000000000000",52264 => "0000000000000000",
52265 => "0000000000000000",52266 => "0000000000000000",
52267 => "0000000000000000",52268 => "0000000000000000",
52269 => "0000000000000000",52270 => "0000000000000000",
52271 => "0000000000000000",52272 => "0000000000000000",
52273 => "0000000000000000",52274 => "0000000000000000",
52275 => "0000000000000000",52276 => "0000000000000000",
52277 => "0000000000000000",52278 => "0000000000000000",
52279 => "0000000000000000",52280 => "0000000000000000",
52281 => "0000000000000000",52282 => "0000000000000000",
52283 => "0000000000000000",52284 => "0000000000000000",
52285 => "0000000000000000",52286 => "0000000000000000",
52287 => "0000000000000000",52288 => "0000000000000000",
52289 => "0000000000000000",52290 => "0000000000000000",
52291 => "0000000000000000",52292 => "0000000000000000",
52293 => "0000000000000000",52294 => "0000000000000000",
52295 => "0000000000000000",52296 => "0000000000000000",
52297 => "0000000000000000",52298 => "0000000000000000",
52299 => "0000000000000000",52300 => "0000000000000000",
52301 => "0000000000000000",52302 => "0000000000000000",
52303 => "0000000000000000",52304 => "0000000000000000",
52305 => "0000000000000000",52306 => "0000000000000000",
52307 => "0000000000000000",52308 => "0000000000000000",
52309 => "0000000000000000",52310 => "0000000000000000",
52311 => "0000000000000000",52312 => "0000000000000000",
52313 => "0000000000000000",52314 => "0000000000000000",
52315 => "0000000000000000",52316 => "0000000000000000",
52317 => "0000000000000000",52318 => "0000000000000000",
52319 => "0000000000000000",52320 => "0000000000000000",
52321 => "0000000000000000",52322 => "0000000000000000",
52323 => "0000000000000000",52324 => "0000000000000000",
52325 => "0000000000000000",52326 => "0000000000000000",
52327 => "0000000000000000",52328 => "0000000000000000",
52329 => "0000000000000000",52330 => "0000000000000000",
52331 => "0000000000000000",52332 => "0000000000000000",
52333 => "0000000000000000",52334 => "0000000000000000",
52335 => "0000000000000000",52336 => "0000000000000000",
52337 => "0000000000000000",52338 => "0000000000000000",
52339 => "0000000000000000",52340 => "0000000000000000",
52341 => "0000000000000000",52342 => "0000000000000000",
52343 => "0000000000000000",52344 => "0000000000000000",
52345 => "0000000000000000",52346 => "0000000000000000",
52347 => "0000000000000000",52348 => "0000000000000000",
52349 => "0000000000000000",52350 => "0000000000000000",
52351 => "0000000000000000",52352 => "0000000000000000",
52353 => "0000000000000000",52354 => "0000000000000000",
52355 => "0000000000000000",52356 => "0000000000000000",
52357 => "0000000000000000",52358 => "0000000000000000",
52359 => "0000000000000000",52360 => "0000000000000000",
52361 => "0000000000000000",52362 => "0000000000000000",
52363 => "0000000000000000",52364 => "0000000000000000",
52365 => "0000000000000000",52366 => "0000000000000000",
52367 => "0000000000000000",52368 => "0000000000000000",
52369 => "0000000000000000",52370 => "0000000000000000",
52371 => "0000000000000000",52372 => "0000000000000000",
52373 => "0000000000000000",52374 => "0000000000000000",
52375 => "0000000000000000",52376 => "0000000000000000",
52377 => "0000000000000000",52378 => "0000000000000000",
52379 => "0000000000000000",52380 => "0000000000000000",
52381 => "0000000000000000",52382 => "0000000000000000",
52383 => "0000000000000000",52384 => "0000000000000000",
52385 => "0000000000000000",52386 => "0000000000000000",
52387 => "0000000000000000",52388 => "0000000000000000",
52389 => "0000000000000000",52390 => "0000000000000000",
52391 => "0000000000000000",52392 => "0000000000000000",
52393 => "0000000000000000",52394 => "0000000000000000",
52395 => "0000000000000000",52396 => "0000000000000000",
52397 => "0000000000000000",52398 => "0000000000000000",
52399 => "0000000000000000",52400 => "0000000000000000",
52401 => "0000000000000000",52402 => "0000000000000000",
52403 => "0000000000000000",52404 => "0000000000000000",
52405 => "0000000000000000",52406 => "0000000000000000",
52407 => "0000000000000000",52408 => "0000000000000000",
52409 => "0000000000000000",52410 => "0000000000000000",
52411 => "0000000000000000",52412 => "0000000000000000",
52413 => "0000000000000000",52414 => "0000000000000000",
52415 => "0000000000000000",52416 => "0000000000000000",
52417 => "0000000000000000",52418 => "0000000000000000",
52419 => "0000000000000000",52420 => "0000000000000000",
52421 => "0000000000000000",52422 => "0000000000000000",
52423 => "0000000000000000",52424 => "0000000000000000",
52425 => "0000000000000000",52426 => "0000000000000000",
52427 => "0000000000000000",52428 => "0000000000000000",
52429 => "0000000000000000",52430 => "0000000000000000",
52431 => "0000000000000000",52432 => "0000000000000000",
52433 => "0000000000000000",52434 => "0000000000000000",
52435 => "0000000000000000",52436 => "0000000000000000",
52437 => "0000000000000000",52438 => "0000000000000000",
52439 => "0000000000000000",52440 => "0000000000000000",
52441 => "0000000000000000",52442 => "0000000000000000",
52443 => "0000000000000000",52444 => "0000000000000000",
52445 => "0000000000000000",52446 => "0000000000000000",
52447 => "0000000000000000",52448 => "0000000000000000",
52449 => "0000000000000000",52450 => "0000000000000000",
52451 => "0000000000000000",52452 => "0000000000000000",
52453 => "0000000000000000",52454 => "0000000000000000",
52455 => "0000000000000000",52456 => "0000000000000000",
52457 => "0000000000000000",52458 => "0000000000000000",
52459 => "0000000000000000",52460 => "0000000000000000",
52461 => "0000000000000000",52462 => "0000000000000000",
52463 => "0000000000000000",52464 => "0000000000000000",
52465 => "0000000000000000",52466 => "0000000000000000",
52467 => "0000000000000000",52468 => "0000000000000000",
52469 => "0000000000000000",52470 => "0000000000000000",
52471 => "0000000000000000",52472 => "0000000000000000",
52473 => "0000000000000000",52474 => "0000000000000000",
52475 => "0000000000000000",52476 => "0000000000000000",
52477 => "0000000000000000",52478 => "0000000000000000",
52479 => "0000000000000000",52480 => "0000000000000000",
52481 => "0000000000000000",52482 => "0000000000000000",
52483 => "0000000000000000",52484 => "0000000000000000",
52485 => "0000000000000000",52486 => "0000000000000000",
52487 => "0000000000000000",52488 => "0000000000000000",
52489 => "0000000000000000",52490 => "0000000000000000",
52491 => "0000000000000000",52492 => "0000000000000000",
52493 => "0000000000000000",52494 => "0000000000000000",
52495 => "0000000000000000",52496 => "0000000000000000",
52497 => "0000000000000000",52498 => "0000000000000000",
52499 => "0000000000000000",52500 => "0000000000000000",
52501 => "0000000000000000",52502 => "0000000000000000",
52503 => "0000000000000000",52504 => "0000000000000000",
52505 => "0000000000000000",52506 => "0000000000000000",
52507 => "0000000000000000",52508 => "0000000000000000",
52509 => "0000000000000000",52510 => "0000000000000000",
52511 => "0000000000000000",52512 => "0000000000000000",
52513 => "0000000000000000",52514 => "0000000000000000",
52515 => "0000000000000000",52516 => "0000000000000000",
52517 => "0000000000000000",52518 => "0000000000000000",
52519 => "0000000000000000",52520 => "0000000000000000",
52521 => "0000000000000000",52522 => "0000000000000000",
52523 => "0000000000000000",52524 => "0000000000000000",
52525 => "0000000000000000",52526 => "0000000000000000",
52527 => "0000000000000000",52528 => "0000000000000000",
52529 => "0000000000000000",52530 => "0000000000000000",
52531 => "0000000000000000",52532 => "0000000000000000",
52533 => "0000000000000000",52534 => "0000000000000000",
52535 => "0000000000000000",52536 => "0000000000000000",
52537 => "0000000000000000",52538 => "0000000000000000",
52539 => "0000000000000000",52540 => "0000000000000000",
52541 => "0000000000000000",52542 => "0000000000000000",
52543 => "0000000000000000",52544 => "0000000000000000",
52545 => "0000000000000000",52546 => "0000000000000000",
52547 => "0000000000000000",52548 => "0000000000000000",
52549 => "0000000000000000",52550 => "0000000000000000",
52551 => "0000000000000000",52552 => "0000000000000000",
52553 => "0000000000000000",52554 => "0000000000000000",
52555 => "0000000000000000",52556 => "0000000000000000",
52557 => "0000000000000000",52558 => "0000000000000000",
52559 => "0000000000000000",52560 => "0000000000000000",
52561 => "0000000000000000",52562 => "0000000000000000",
52563 => "0000000000000000",52564 => "0000000000000000",
52565 => "0000000000000000",52566 => "0000000000000000",
52567 => "0000000000000000",52568 => "0000000000000000",
52569 => "0000000000000000",52570 => "0000000000000000",
52571 => "0000000000000000",52572 => "0000000000000000",
52573 => "0000000000000000",52574 => "0000000000000000",
52575 => "0000000000000000",52576 => "0000000000000000",
52577 => "0000000000000000",52578 => "0000000000000000",
52579 => "0000000000000000",52580 => "0000000000000000",
52581 => "0000000000000000",52582 => "0000000000000000",
52583 => "0000000000000000",52584 => "0000000000000000",
52585 => "0000000000000000",52586 => "0000000000000000",
52587 => "0000000000000000",52588 => "0000000000000000",
52589 => "0000000000000000",52590 => "0000000000000000",
52591 => "0000000000000000",52592 => "0000000000000000",
52593 => "0000000000000000",52594 => "0000000000000000",
52595 => "0000000000000000",52596 => "0000000000000000",
52597 => "0000000000000000",52598 => "0000000000000000",
52599 => "0000000000000000",52600 => "0000000000000000",
52601 => "0000000000000000",52602 => "0000000000000000",
52603 => "0000000000000000",52604 => "0000000000000000",
52605 => "0000000000000000",52606 => "0000000000000000",
52607 => "0000000000000000",52608 => "0000000000000000",
52609 => "0000000000000000",52610 => "0000000000000000",
52611 => "0000000000000000",52612 => "0000000000000000",
52613 => "0000000000000000",52614 => "0000000000000000",
52615 => "0000000000000000",52616 => "0000000000000000",
52617 => "0000000000000000",52618 => "0000000000000000",
52619 => "0000000000000000",52620 => "0000000000000000",
52621 => "0000000000000000",52622 => "0000000000000000",
52623 => "0000000000000000",52624 => "0000000000000000",
52625 => "0000000000000000",52626 => "0000000000000000",
52627 => "0000000000000000",52628 => "0000000000000000",
52629 => "0000000000000000",52630 => "0000000000000000",
52631 => "0000000000000000",52632 => "0000000000000000",
52633 => "0000000000000000",52634 => "0000000000000000",
52635 => "0000000000000000",52636 => "0000000000000000",
52637 => "0000000000000000",52638 => "0000000000000000",
52639 => "0000000000000000",52640 => "0000000000000000",
52641 => "0000000000000000",52642 => "0000000000000000",
52643 => "0000000000000000",52644 => "0000000000000000",
52645 => "0000000000000000",52646 => "0000000000000000",
52647 => "0000000000000000",52648 => "0000000000000000",
52649 => "0000000000000000",52650 => "0000000000000000",
52651 => "0000000000000000",52652 => "0000000000000000",
52653 => "0000000000000000",52654 => "0000000000000000",
52655 => "0000000000000000",52656 => "0000000000000000",
52657 => "0000000000000000",52658 => "0000000000000000",
52659 => "0000000000000000",52660 => "0000000000000000",
52661 => "0000000000000000",52662 => "0000000000000000",
52663 => "0000000000000000",52664 => "0000000000000000",
52665 => "0000000000000000",52666 => "0000000000000000",
52667 => "0000000000000000",52668 => "0000000000000000",
52669 => "0000000000000000",52670 => "0000000000000000",
52671 => "0000000000000000",52672 => "0000000000000000",
52673 => "0000000000000000",52674 => "0000000000000000",
52675 => "0000000000000000",52676 => "0000000000000000",
52677 => "0000000000000000",52678 => "0000000000000000",
52679 => "0000000000000000",52680 => "0000000000000000",
52681 => "0000000000000000",52682 => "0000000000000000",
52683 => "0000000000000000",52684 => "0000000000000000",
52685 => "0000000000000000",52686 => "0000000000000000",
52687 => "0000000000000000",52688 => "0000000000000000",
52689 => "0000000000000000",52690 => "0000000000000000",
52691 => "0000000000000000",52692 => "0000000000000000",
52693 => "0000000000000000",52694 => "0000000000000000",
52695 => "0000000000000000",52696 => "0000000000000000",
52697 => "0000000000000000",52698 => "0000000000000000",
52699 => "0000000000000000",52700 => "0000000000000000",
52701 => "0000000000000000",52702 => "0000000000000000",
52703 => "0000000000000000",52704 => "0000000000000000",
52705 => "0000000000000000",52706 => "0000000000000000",
52707 => "0000000000000000",52708 => "0000000000000000",
52709 => "0000000000000000",52710 => "0000000000000000",
52711 => "0000000000000000",52712 => "0000000000000000",
52713 => "0000000000000000",52714 => "0000000000000000",
52715 => "0000000000000000",52716 => "0000000000000000",
52717 => "0000000000000000",52718 => "0000000000000000",
52719 => "0000000000000000",52720 => "0000000000000000",
52721 => "0000000000000000",52722 => "0000000000000000",
52723 => "0000000000000000",52724 => "0000000000000000",
52725 => "0000000000000000",52726 => "0000000000000000",
52727 => "0000000000000000",52728 => "0000000000000000",
52729 => "0000000000000000",52730 => "0000000000000000",
52731 => "0000000000000000",52732 => "0000000000000000",
52733 => "0000000000000000",52734 => "0000000000000000",
52735 => "0000000000000000",52736 => "0000000000000000",
52737 => "0000000000000000",52738 => "0000000000000000",
52739 => "0000000000000000",52740 => "0000000000000000",
52741 => "0000000000000000",52742 => "0000000000000000",
52743 => "0000000000000000",52744 => "0000000000000000",
52745 => "0000000000000000",52746 => "0000000000000000",
52747 => "0000000000000000",52748 => "0000000000000000",
52749 => "0000000000000000",52750 => "0000000000000000",
52751 => "0000000000000000",52752 => "0000000000000000",
52753 => "0000000000000000",52754 => "0000000000000000",
52755 => "0000000000000000",52756 => "0000000000000000",
52757 => "0000000000000000",52758 => "0000000000000000",
52759 => "0000000000000000",52760 => "0000000000000000",
52761 => "0000000000000000",52762 => "0000000000000000",
52763 => "0000000000000000",52764 => "0000000000000000",
52765 => "0000000000000000",52766 => "0000000000000000",
52767 => "0000000000000000",52768 => "0000000000000000",
52769 => "0000000000000000",52770 => "0000000000000000",
52771 => "0000000000000000",52772 => "0000000000000000",
52773 => "0000000000000000",52774 => "0000000000000000",
52775 => "0000000000000000",52776 => "0000000000000000",
52777 => "0000000000000000",52778 => "0000000000000000",
52779 => "0000000000000000",52780 => "0000000000000000",
52781 => "0000000000000000",52782 => "0000000000000000",
52783 => "0000000000000000",52784 => "0000000000000000",
52785 => "0000000000000000",52786 => "0000000000000000",
52787 => "0000000000000000",52788 => "0000000000000000",
52789 => "0000000000000000",52790 => "0000000000000000",
52791 => "0000000000000000",52792 => "0000000000000000",
52793 => "0000000000000000",52794 => "0000000000000000",
52795 => "0000000000000000",52796 => "0000000000000000",
52797 => "0000000000000000",52798 => "0000000000000000",
52799 => "0000000000000000",52800 => "0000000000000000",
52801 => "0000000000000000",52802 => "0000000000000000",
52803 => "0000000000000000",52804 => "0000000000000000",
52805 => "0000000000000000",52806 => "0000000000000000",
52807 => "0000000000000000",52808 => "0000000000000000",
52809 => "0000000000000000",52810 => "0000000000000000",
52811 => "0000000000000000",52812 => "0000000000000000",
52813 => "0000000000000000",52814 => "0000000000000000",
52815 => "0000000000000000",52816 => "0000000000000000",
52817 => "0000000000000000",52818 => "0000000000000000",
52819 => "0000000000000000",52820 => "0000000000000000",
52821 => "0000000000000000",52822 => "0000000000000000",
52823 => "0000000000000000",52824 => "0000000000000000",
52825 => "0000000000000000",52826 => "0000000000000000",
52827 => "0000000000000000",52828 => "0000000000000000",
52829 => "0000000000000000",52830 => "0000000000000000",
52831 => "0000000000000000",52832 => "0000000000000000",
52833 => "0000000000000000",52834 => "0000000000000000",
52835 => "0000000000000000",52836 => "0000000000000000",
52837 => "0000000000000000",52838 => "0000000000000000",
52839 => "0000000000000000",52840 => "0000000000000000",
52841 => "0000000000000000",52842 => "0000000000000000",
52843 => "0000000000000000",52844 => "0000000000000000",
52845 => "0000000000000000",52846 => "0000000000000000",
52847 => "0000000000000000",52848 => "0000000000000000",
52849 => "0000000000000000",52850 => "0000000000000000",
52851 => "0000000000000000",52852 => "0000000000000000",
52853 => "0000000000000000",52854 => "0000000000000000",
52855 => "0000000000000000",52856 => "0000000000000000",
52857 => "0000000000000000",52858 => "0000000000000000",
52859 => "0000000000000000",52860 => "0000000000000000",
52861 => "0000000000000000",52862 => "0000000000000000",
52863 => "0000000000000000",52864 => "0000000000000000",
52865 => "0000000000000000",52866 => "0000000000000000",
52867 => "0000000000000000",52868 => "0000000000000000",
52869 => "0000000000000000",52870 => "0000000000000000",
52871 => "0000000000000000",52872 => "0000000000000000",
52873 => "0000000000000000",52874 => "0000000000000000",
52875 => "0000000000000000",52876 => "0000000000000000",
52877 => "0000000000000000",52878 => "0000000000000000",
52879 => "0000000000000000",52880 => "0000000000000000",
52881 => "0000000000000000",52882 => "0000000000000000",
52883 => "0000000000000000",52884 => "0000000000000000",
52885 => "0000000000000000",52886 => "0000000000000000",
52887 => "0000000000000000",52888 => "0000000000000000",
52889 => "0000000000000000",52890 => "0000000000000000",
52891 => "0000000000000000",52892 => "0000000000000000",
52893 => "0000000000000000",52894 => "0000000000000000",
52895 => "0000000000000000",52896 => "0000000000000000",
52897 => "0000000000000000",52898 => "0000000000000000",
52899 => "0000000000000000",52900 => "0000000000000000",
52901 => "0000000000000000",52902 => "0000000000000000",
52903 => "0000000000000000",52904 => "0000000000000000",
52905 => "0000000000000000",52906 => "0000000000000000",
52907 => "0000000000000000",52908 => "0000000000000000",
52909 => "0000000000000000",52910 => "0000000000000000",
52911 => "0000000000000000",52912 => "0000000000000000",
52913 => "0000000000000000",52914 => "0000000000000000",
52915 => "0000000000000000",52916 => "0000000000000000",
52917 => "0000000000000000",52918 => "0000000000000000",
52919 => "0000000000000000",52920 => "0000000000000000",
52921 => "0000000000000000",52922 => "0000000000000000",
52923 => "0000000000000000",52924 => "0000000000000000",
52925 => "0000000000000000",52926 => "0000000000000000",
52927 => "0000000000000000",52928 => "0000000000000000",
52929 => "0000000000000000",52930 => "0000000000000000",
52931 => "0000000000000000",52932 => "0000000000000000",
52933 => "0000000000000000",52934 => "0000000000000000",
52935 => "0000000000000000",52936 => "0000000000000000",
52937 => "0000000000000000",52938 => "0000000000000000",
52939 => "0000000000000000",52940 => "0000000000000000",
52941 => "0000000000000000",52942 => "0000000000000000",
52943 => "0000000000000000",52944 => "0000000000000000",
52945 => "0000000000000000",52946 => "0000000000000000",
52947 => "0000000000000000",52948 => "0000000000000000",
52949 => "0000000000000000",52950 => "0000000000000000",
52951 => "0000000000000000",52952 => "0000000000000000",
52953 => "0000000000000000",52954 => "0000000000000000",
52955 => "0000000000000000",52956 => "0000000000000000",
52957 => "0000000000000000",52958 => "0000000000000000",
52959 => "0000000000000000",52960 => "0000000000000000",
52961 => "0000000000000000",52962 => "0000000000000000",
52963 => "0000000000000000",52964 => "0000000000000000",
52965 => "0000000000000000",52966 => "0000000000000000",
52967 => "0000000000000000",52968 => "0000000000000000",
52969 => "0000000000000000",52970 => "0000000000000000",
52971 => "0000000000000000",52972 => "0000000000000000",
52973 => "0000000000000000",52974 => "0000000000000000",
52975 => "0000000000000000",52976 => "0000000000000000",
52977 => "0000000000000000",52978 => "0000000000000000",
52979 => "0000000000000000",52980 => "0000000000000000",
52981 => "0000000000000000",52982 => "0000000000000000",
52983 => "0000000000000000",52984 => "0000000000000000",
52985 => "0000000000000000",52986 => "0000000000000000",
52987 => "0000000000000000",52988 => "0000000000000000",
52989 => "0000000000000000",52990 => "0000000000000000",
52991 => "0000000000000000",52992 => "0000000000000000",
52993 => "0000000000000000",52994 => "0000000000000000",
52995 => "0000000000000000",52996 => "0000000000000000",
52997 => "0000000000000000",52998 => "0000000000000000",
52999 => "0000000000000000",53000 => "0000000000000000",
53001 => "0000000000000000",53002 => "0000000000000000",
53003 => "0000000000000000",53004 => "0000000000000000",
53005 => "0000000000000000",53006 => "0000000000000000",
53007 => "0000000000000000",53008 => "0000000000000000",
53009 => "0000000000000000",53010 => "0000000000000000",
53011 => "0000000000000000",53012 => "0000000000000000",
53013 => "0000000000000000",53014 => "0000000000000000",
53015 => "0000000000000000",53016 => "0000000000000000",
53017 => "0000000000000000",53018 => "0000000000000000",
53019 => "0000000000000000",53020 => "0000000000000000",
53021 => "0000000000000000",53022 => "0000000000000000",
53023 => "0000000000000000",53024 => "0000000000000000",
53025 => "0000000000000000",53026 => "0000000000000000",
53027 => "0000000000000000",53028 => "0000000000000000",
53029 => "0000000000000000",53030 => "0000000000000000",
53031 => "0000000000000000",53032 => "0000000000000000",
53033 => "0000000000000000",53034 => "0000000000000000",
53035 => "0000000000000000",53036 => "0000000000000000",
53037 => "0000000000000000",53038 => "0000000000000000",
53039 => "0000000000000000",53040 => "0000000000000000",
53041 => "0000000000000000",53042 => "0000000000000000",
53043 => "0000000000000000",53044 => "0000000000000000",
53045 => "0000000000000000",53046 => "0000000000000000",
53047 => "0000000000000000",53048 => "0000000000000000",
53049 => "0000000000000000",53050 => "0000000000000000",
53051 => "0000000000000000",53052 => "0000000000000000",
53053 => "0000000000000000",53054 => "0000000000000000",
53055 => "0000000000000000",53056 => "0000000000000000",
53057 => "0000000000000000",53058 => "0000000000000000",
53059 => "0000000000000000",53060 => "0000000000000000",
53061 => "0000000000000000",53062 => "0000000000000000",
53063 => "0000000000000000",53064 => "0000000000000000",
53065 => "0000000000000000",53066 => "0000000000000000",
53067 => "0000000000000000",53068 => "0000000000000000",
53069 => "0000000000000000",53070 => "0000000000000000",
53071 => "0000000000000000",53072 => "0000000000000000",
53073 => "0000000000000000",53074 => "0000000000000000",
53075 => "0000000000000000",53076 => "0000000000000000",
53077 => "0000000000000000",53078 => "0000000000000000",
53079 => "0000000000000000",53080 => "0000000000000000",
53081 => "0000000000000000",53082 => "0000000000000000",
53083 => "0000000000000000",53084 => "0000000000000000",
53085 => "0000000000000000",53086 => "0000000000000000",
53087 => "0000000000000000",53088 => "0000000000000000",
53089 => "0000000000000000",53090 => "0000000000000000",
53091 => "0000000000000000",53092 => "0000000000000000",
53093 => "0000000000000000",53094 => "0000000000000000",
53095 => "0000000000000000",53096 => "0000000000000000",
53097 => "0000000000000000",53098 => "0000000000000000",
53099 => "0000000000000000",53100 => "0000000000000000",
53101 => "0000000000000000",53102 => "0000000000000000",
53103 => "0000000000000000",53104 => "0000000000000000",
53105 => "0000000000000000",53106 => "0000000000000000",
53107 => "0000000000000000",53108 => "0000000000000000",
53109 => "0000000000000000",53110 => "0000000000000000",
53111 => "0000000000000000",53112 => "0000000000000000",
53113 => "0000000000000000",53114 => "0000000000000000",
53115 => "0000000000000000",53116 => "0000000000000000",
53117 => "0000000000000000",53118 => "0000000000000000",
53119 => "0000000000000000",53120 => "0000000000000000",
53121 => "0000000000000000",53122 => "0000000000000000",
53123 => "0000000000000000",53124 => "0000000000000000",
53125 => "0000000000000000",53126 => "0000000000000000",
53127 => "0000000000000000",53128 => "0000000000000000",
53129 => "0000000000000000",53130 => "0000000000000000",
53131 => "0000000000000000",53132 => "0000000000000000",
53133 => "0000000000000000",53134 => "0000000000000000",
53135 => "0000000000000000",53136 => "0000000000000000",
53137 => "0000000000000000",53138 => "0000000000000000",
53139 => "0000000000000000",53140 => "0000000000000000",
53141 => "0000000000000000",53142 => "0000000000000000",
53143 => "0000000000000000",53144 => "0000000000000000",
53145 => "0000000000000000",53146 => "0000000000000000",
53147 => "0000000000000000",53148 => "0000000000000000",
53149 => "0000000000000000",53150 => "0000000000000000",
53151 => "0000000000000000",53152 => "0000000000000000",
53153 => "0000000000000000",53154 => "0000000000000000",
53155 => "0000000000000000",53156 => "0000000000000000",
53157 => "0000000000000000",53158 => "0000000000000000",
53159 => "0000000000000000",53160 => "0000000000000000",
53161 => "0000000000000000",53162 => "0000000000000000",
53163 => "0000000000000000",53164 => "0000000000000000",
53165 => "0000000000000000",53166 => "0000000000000000",
53167 => "0000000000000000",53168 => "0000000000000000",
53169 => "0000000000000000",53170 => "0000000000000000",
53171 => "0000000000000000",53172 => "0000000000000000",
53173 => "0000000000000000",53174 => "0000000000000000",
53175 => "0000000000000000",53176 => "0000000000000000",
53177 => "0000000000000000",53178 => "0000000000000000",
53179 => "0000000000000000",53180 => "0000000000000000",
53181 => "0000000000000000",53182 => "0000000000000000",
53183 => "0000000000000000",53184 => "0000000000000000",
53185 => "0000000000000000",53186 => "0000000000000000",
53187 => "0000000000000000",53188 => "0000000000000000",
53189 => "0000000000000000",53190 => "0000000000000000",
53191 => "0000000000000000",53192 => "0000000000000000",
53193 => "0000000000000000",53194 => "0000000000000000",
53195 => "0000000000000000",53196 => "0000000000000000",
53197 => "0000000000000000",53198 => "0000000000000000",
53199 => "0000000000000000",53200 => "0000000000000000",
53201 => "0000000000000000",53202 => "0000000000000000",
53203 => "0000000000000000",53204 => "0000000000000000",
53205 => "0000000000000000",53206 => "0000000000000000",
53207 => "0000000000000000",53208 => "0000000000000000",
53209 => "0000000000000000",53210 => "0000000000000000",
53211 => "0000000000000000",53212 => "0000000000000000",
53213 => "0000000000000000",53214 => "0000000000000000",
53215 => "0000000000000000",53216 => "0000000000000000",
53217 => "0000000000000000",53218 => "0000000000000000",
53219 => "0000000000000000",53220 => "0000000000000000",
53221 => "0000000000000000",53222 => "0000000000000000",
53223 => "0000000000000000",53224 => "0000000000000000",
53225 => "0000000000000000",53226 => "0000000000000000",
53227 => "0000000000000000",53228 => "0000000000000000",
53229 => "0000000000000000",53230 => "0000000000000000",
53231 => "0000000000000000",53232 => "0000000000000000",
53233 => "0000000000000000",53234 => "0000000000000000",
53235 => "0000000000000000",53236 => "0000000000000000",
53237 => "0000000000000000",53238 => "0000000000000000",
53239 => "0000000000000000",53240 => "0000000000000000",
53241 => "0000000000000000",53242 => "0000000000000000",
53243 => "0000000000000000",53244 => "0000000000000000",
53245 => "0000000000000000",53246 => "0000000000000000",
53247 => "0000000000000000",53248 => "0000000000000000",
53249 => "0000000000000000",53250 => "0000000000000000",
53251 => "0000000000000000",53252 => "0000000000000000",
53253 => "0000000000000000",53254 => "0000000000000000",
53255 => "0000000000000000",53256 => "0000000000000000",
53257 => "0000000000000000",53258 => "0000000000000000",
53259 => "0000000000000000",53260 => "0000000000000000",
53261 => "0000000000000000",53262 => "0000000000000000",
53263 => "0000000000000000",53264 => "0000000000000000",
53265 => "0000000000000000",53266 => "0000000000000000",
53267 => "0000000000000000",53268 => "0000000000000000",
53269 => "0000000000000000",53270 => "0000000000000000",
53271 => "0000000000000000",53272 => "0000000000000000",
53273 => "0000000000000000",53274 => "0000000000000000",
53275 => "0000000000000000",53276 => "0000000000000000",
53277 => "0000000000000000",53278 => "0000000000000000",
53279 => "0000000000000000",53280 => "0000000000000000",
53281 => "0000000000000000",53282 => "0000000000000000",
53283 => "0000000000000000",53284 => "0000000000000000",
53285 => "0000000000000000",53286 => "0000000000000000",
53287 => "0000000000000000",53288 => "0000000000000000",
53289 => "0000000000000000",53290 => "0000000000000000",
53291 => "0000000000000000",53292 => "0000000000000000",
53293 => "0000000000000000",53294 => "0000000000000000",
53295 => "0000000000000000",53296 => "0000000000000000",
53297 => "0000000000000000",53298 => "0000000000000000",
53299 => "0000000000000000",53300 => "0000000000000000",
53301 => "0000000000000000",53302 => "0000000000000000",
53303 => "0000000000000000",53304 => "0000000000000000",
53305 => "0000000000000000",53306 => "0000000000000000",
53307 => "0000000000000000",53308 => "0000000000000000",
53309 => "0000000000000000",53310 => "0000000000000000",
53311 => "0000000000000000",53312 => "0000000000000000",
53313 => "0000000000000000",53314 => "0000000000000000",
53315 => "0000000000000000",53316 => "0000000000000000",
53317 => "0000000000000000",53318 => "0000000000000000",
53319 => "0000000000000000",53320 => "0000000000000000",
53321 => "0000000000000000",53322 => "0000000000000000",
53323 => "0000000000000000",53324 => "0000000000000000",
53325 => "0000000000000000",53326 => "0000000000000000",
53327 => "0000000000000000",53328 => "0000000000000000",
53329 => "0000000000000000",53330 => "0000000000000000",
53331 => "0000000000000000",53332 => "0000000000000000",
53333 => "0000000000000000",53334 => "0000000000000000",
53335 => "0000000000000000",53336 => "0000000000000000",
53337 => "0000000000000000",53338 => "0000000000000000",
53339 => "0000000000000000",53340 => "0000000000000000",
53341 => "0000000000000000",53342 => "0000000000000000",
53343 => "0000000000000000",53344 => "0000000000000000",
53345 => "0000000000000000",53346 => "0000000000000000",
53347 => "0000000000000000",53348 => "0000000000000000",
53349 => "0000000000000000",53350 => "0000000000000000",
53351 => "0000000000000000",53352 => "0000000000000000",
53353 => "0000000000000000",53354 => "0000000000000000",
53355 => "0000000000000000",53356 => "0000000000000000",
53357 => "0000000000000000",53358 => "0000000000000000",
53359 => "0000000000000000",53360 => "0000000000000000",
53361 => "0000000000000000",53362 => "0000000000000000",
53363 => "0000000000000000",53364 => "0000000000000000",
53365 => "0000000000000000",53366 => "0000000000000000",
53367 => "0000000000000000",53368 => "0000000000000000",
53369 => "0000000000000000",53370 => "0000000000000000",
53371 => "0000000000000000",53372 => "0000000000000000",
53373 => "0000000000000000",53374 => "0000000000000000",
53375 => "0000000000000000",53376 => "0000000000000000",
53377 => "0000000000000000",53378 => "0000000000000000",
53379 => "0000000000000000",53380 => "0000000000000000",
53381 => "0000000000000000",53382 => "0000000000000000",
53383 => "0000000000000000",53384 => "0000000000000000",
53385 => "0000000000000000",53386 => "0000000000000000",
53387 => "0000000000000000",53388 => "0000000000000000",
53389 => "0000000000000000",53390 => "0000000000000000",
53391 => "0000000000000000",53392 => "0000000000000000",
53393 => "0000000000000000",53394 => "0000000000000000",
53395 => "0000000000000000",53396 => "0000000000000000",
53397 => "0000000000000000",53398 => "0000000000000000",
53399 => "0000000000000000",53400 => "0000000000000000",
53401 => "0000000000000000",53402 => "0000000000000000",
53403 => "0000000000000000",53404 => "0000000000000000",
53405 => "0000000000000000",53406 => "0000000000000000",
53407 => "0000000000000000",53408 => "0000000000000000",
53409 => "0000000000000000",53410 => "0000000000000000",
53411 => "0000000000000000",53412 => "0000000000000000",
53413 => "0000000000000000",53414 => "0000000000000000",
53415 => "0000000000000000",53416 => "0000000000000000",
53417 => "0000000000000000",53418 => "0000000000000000",
53419 => "0000000000000000",53420 => "0000000000000000",
53421 => "0000000000000000",53422 => "0000000000000000",
53423 => "0000000000000000",53424 => "0000000000000000",
53425 => "0000000000000000",53426 => "0000000000000000",
53427 => "0000000000000000",53428 => "0000000000000000",
53429 => "0000000000000000",53430 => "0000000000000000",
53431 => "0000000000000000",53432 => "0000000000000000",
53433 => "0000000000000000",53434 => "0000000000000000",
53435 => "0000000000000000",53436 => "0000000000000000",
53437 => "0000000000000000",53438 => "0000000000000000",
53439 => "0000000000000000",53440 => "0000000000000000",
53441 => "0000000000000000",53442 => "0000000000000000",
53443 => "0000000000000000",53444 => "0000000000000000",
53445 => "0000000000000000",53446 => "0000000000000000",
53447 => "0000000000000000",53448 => "0000000000000000",
53449 => "0000000000000000",53450 => "0000000000000000",
53451 => "0000000000000000",53452 => "0000000000000000",
53453 => "0000000000000000",53454 => "0000000000000000",
53455 => "0000000000000000",53456 => "0000000000000000",
53457 => "0000000000000000",53458 => "0000000000000000",
53459 => "0000000000000000",53460 => "0000000000000000",
53461 => "0000000000000000",53462 => "0000000000000000",
53463 => "0000000000000000",53464 => "0000000000000000",
53465 => "0000000000000000",53466 => "0000000000000000",
53467 => "0000000000000000",53468 => "0000000000000000",
53469 => "0000000000000000",53470 => "0000000000000000",
53471 => "0000000000000000",53472 => "0000000000000000",
53473 => "0000000000000000",53474 => "0000000000000000",
53475 => "0000000000000000",53476 => "0000000000000000",
53477 => "0000000000000000",53478 => "0000000000000000",
53479 => "0000000000000000",53480 => "0000000000000000",
53481 => "0000000000000000",53482 => "0000000000000000",
53483 => "0000000000000000",53484 => "0000000000000000",
53485 => "0000000000000000",53486 => "0000000000000000",
53487 => "0000000000000000",53488 => "0000000000000000",
53489 => "0000000000000000",53490 => "0000000000000000",
53491 => "0000000000000000",53492 => "0000000000000000",
53493 => "0000000000000000",53494 => "0000000000000000",
53495 => "0000000000000000",53496 => "0000000000000000",
53497 => "0000000000000000",53498 => "0000000000000000",
53499 => "0000000000000000",53500 => "0000000000000000",
53501 => "0000000000000000",53502 => "0000000000000000",
53503 => "0000000000000000",53504 => "0000000000000000",
53505 => "0000000000000000",53506 => "0000000000000000",
53507 => "0000000000000000",53508 => "0000000000000000",
53509 => "0000000000000000",53510 => "0000000000000000",
53511 => "0000000000000000",53512 => "0000000000000000",
53513 => "0000000000000000",53514 => "0000000000000000",
53515 => "0000000000000000",53516 => "0000000000000000",
53517 => "0000000000000000",53518 => "0000000000000000",
53519 => "0000000000000000",53520 => "0000000000000000",
53521 => "0000000000000000",53522 => "0000000000000000",
53523 => "0000000000000000",53524 => "0000000000000000",
53525 => "0000000000000000",53526 => "0000000000000000",
53527 => "0000000000000000",53528 => "0000000000000000",
53529 => "0000000000000000",53530 => "0000000000000000",
53531 => "0000000000000000",53532 => "0000000000000000",
53533 => "0000000000000000",53534 => "0000000000000000",
53535 => "0000000000000000",53536 => "0000000000000000",
53537 => "0000000000000000",53538 => "0000000000000000",
53539 => "0000000000000000",53540 => "0000000000000000",
53541 => "0000000000000000",53542 => "0000000000000000",
53543 => "0000000000000000",53544 => "0000000000000000",
53545 => "0000000000000000",53546 => "0000000000000000",
53547 => "0000000000000000",53548 => "0000000000000000",
53549 => "0000000000000000",53550 => "0000000000000000",
53551 => "0000000000000000",53552 => "0000000000000000",
53553 => "0000000000000000",53554 => "0000000000000000",
53555 => "0000000000000000",53556 => "0000000000000000",
53557 => "0000000000000000",53558 => "0000000000000000",
53559 => "0000000000000000",53560 => "0000000000000000",
53561 => "0000000000000000",53562 => "0000000000000000",
53563 => "0000000000000000",53564 => "0000000000000000",
53565 => "0000000000000000",53566 => "0000000000000000",
53567 => "0000000000000000",53568 => "0000000000000000",
53569 => "0000000000000000",53570 => "0000000000000000",
53571 => "0000000000000000",53572 => "0000000000000000",
53573 => "0000000000000000",53574 => "0000000000000000",
53575 => "0000000000000000",53576 => "0000000000000000",
53577 => "0000000000000000",53578 => "0000000000000000",
53579 => "0000000000000000",53580 => "0000000000000000",
53581 => "0000000000000000",53582 => "0000000000000000",
53583 => "0000000000000000",53584 => "0000000000000000",
53585 => "0000000000000000",53586 => "0000000000000000",
53587 => "0000000000000000",53588 => "0000000000000000",
53589 => "0000000000000000",53590 => "0000000000000000",
53591 => "0000000000000000",53592 => "0000000000000000",
53593 => "0000000000000000",53594 => "0000000000000000",
53595 => "0000000000000000",53596 => "0000000000000000",
53597 => "0000000000000000",53598 => "0000000000000000",
53599 => "0000000000000000",53600 => "0000000000000000",
53601 => "0000000000000000",53602 => "0000000000000000",
53603 => "0000000000000000",53604 => "0000000000000000",
53605 => "0000000000000000",53606 => "0000000000000000",
53607 => "0000000000000000",53608 => "0000000000000000",
53609 => "0000000000000000",53610 => "0000000000000000",
53611 => "0000000000000000",53612 => "0000000000000000",
53613 => "0000000000000000",53614 => "0000000000000000",
53615 => "0000000000000000",53616 => "0000000000000000",
53617 => "0000000000000000",53618 => "0000000000000000",
53619 => "0000000000000000",53620 => "0000000000000000",
53621 => "0000000000000000",53622 => "0000000000000000",
53623 => "0000000000000000",53624 => "0000000000000000",
53625 => "0000000000000000",53626 => "0000000000000000",
53627 => "0000000000000000",53628 => "0000000000000000",
53629 => "0000000000000000",53630 => "0000000000000000",
53631 => "0000000000000000",53632 => "0000000000000000",
53633 => "0000000000000000",53634 => "0000000000000000",
53635 => "0000000000000000",53636 => "0000000000000000",
53637 => "0000000000000000",53638 => "0000000000000000",
53639 => "0000000000000000",53640 => "0000000000000000",
53641 => "0000000000000000",53642 => "0000000000000000",
53643 => "0000000000000000",53644 => "0000000000000000",
53645 => "0000000000000000",53646 => "0000000000000000",
53647 => "0000000000000000",53648 => "0000000000000000",
53649 => "0000000000000000",53650 => "0000000000000000",
53651 => "0000000000000000",53652 => "0000000000000000",
53653 => "0000000000000000",53654 => "0000000000000000",
53655 => "0000000000000000",53656 => "0000000000000000",
53657 => "0000000000000000",53658 => "0000000000000000",
53659 => "0000000000000000",53660 => "0000000000000000",
53661 => "0000000000000000",53662 => "0000000000000000",
53663 => "0000000000000000",53664 => "0000000000000000",
53665 => "0000000000000000",53666 => "0000000000000000",
53667 => "0000000000000000",53668 => "0000000000000000",
53669 => "0000000000000000",53670 => "0000000000000000",
53671 => "0000000000000000",53672 => "0000000000000000",
53673 => "0000000000000000",53674 => "0000000000000000",
53675 => "0000000000000000",53676 => "0000000000000000",
53677 => "0000000000000000",53678 => "0000000000000000",
53679 => "0000000000000000",53680 => "0000000000000000",
53681 => "0000000000000000",53682 => "0000000000000000",
53683 => "0000000000000000",53684 => "0000000000000000",
53685 => "0000000000000000",53686 => "0000000000000000",
53687 => "0000000000000000",53688 => "0000000000000000",
53689 => "0000000000000000",53690 => "0000000000000000",
53691 => "0000000000000000",53692 => "0000000000000000",
53693 => "0000000000000000",53694 => "0000000000000000",
53695 => "0000000000000000",53696 => "0000000000000000",
53697 => "0000000000000000",53698 => "0000000000000000",
53699 => "0000000000000000",53700 => "0000000000000000",
53701 => "0000000000000000",53702 => "0000000000000000",
53703 => "0000000000000000",53704 => "0000000000000000",
53705 => "0000000000000000",53706 => "0000000000000000",
53707 => "0000000000000000",53708 => "0000000000000000",
53709 => "0000000000000000",53710 => "0000000000000000",
53711 => "0000000000000000",53712 => "0000000000000000",
53713 => "0000000000000000",53714 => "0000000000000000",
53715 => "0000000000000000",53716 => "0000000000000000",
53717 => "0000000000000000",53718 => "0000000000000000",
53719 => "0000000000000000",53720 => "0000000000000000",
53721 => "0000000000000000",53722 => "0000000000000000",
53723 => "0000000000000000",53724 => "0000000000000000",
53725 => "0000000000000000",53726 => "0000000000000000",
53727 => "0000000000000000",53728 => "0000000000000000",
53729 => "0000000000000000",53730 => "0000000000000000",
53731 => "0000000000000000",53732 => "0000000000000000",
53733 => "0000000000000000",53734 => "0000000000000000",
53735 => "0000000000000000",53736 => "0000000000000000",
53737 => "0000000000000000",53738 => "0000000000000000",
53739 => "0000000000000000",53740 => "0000000000000000",
53741 => "0000000000000000",53742 => "0000000000000000",
53743 => "0000000000000000",53744 => "0000000000000000",
53745 => "0000000000000000",53746 => "0000000000000000",
53747 => "0000000000000000",53748 => "0000000000000000",
53749 => "0000000000000000",53750 => "0000000000000000",
53751 => "0000000000000000",53752 => "0000000000000000",
53753 => "0000000000000000",53754 => "0000000000000000",
53755 => "0000000000000000",53756 => "0000000000000000",
53757 => "0000000000000000",53758 => "0000000000000000",
53759 => "0000000000000000",53760 => "0000000000000000",
53761 => "0000000000000000",53762 => "0000000000000000",
53763 => "0000000000000000",53764 => "0000000000000000",
53765 => "0000000000000000",53766 => "0000000000000000",
53767 => "0000000000000000",53768 => "0000000000000000",
53769 => "0000000000000000",53770 => "0000000000000000",
53771 => "0000000000000000",53772 => "0000000000000000",
53773 => "0000000000000000",53774 => "0000000000000000",
53775 => "0000000000000000",53776 => "0000000000000000",
53777 => "0000000000000000",53778 => "0000000000000000",
53779 => "0000000000000000",53780 => "0000000000000000",
53781 => "0000000000000000",53782 => "0000000000000000",
53783 => "0000000000000000",53784 => "0000000000000000",
53785 => "0000000000000000",53786 => "0000000000000000",
53787 => "0000000000000000",53788 => "0000000000000000",
53789 => "0000000000000000",53790 => "0000000000000000",
53791 => "0000000000000000",53792 => "0000000000000000",
53793 => "0000000000000000",53794 => "0000000000000000",
53795 => "0000000000000000",53796 => "0000000000000000",
53797 => "0000000000000000",53798 => "0000000000000000",
53799 => "0000000000000000",53800 => "0000000000000000",
53801 => "0000000000000000",53802 => "0000000000000000",
53803 => "0000000000000000",53804 => "0000000000000000",
53805 => "0000000000000000",53806 => "0000000000000000",
53807 => "0000000000000000",53808 => "0000000000000000",
53809 => "0000000000000000",53810 => "0000000000000000",
53811 => "0000000000000000",53812 => "0000000000000000",
53813 => "0000000000000000",53814 => "0000000000000000",
53815 => "0000000000000000",53816 => "0000000000000000",
53817 => "0000000000000000",53818 => "0000000000000000",
53819 => "0000000000000000",53820 => "0000000000000000",
53821 => "0000000000000000",53822 => "0000000000000000",
53823 => "0000000000000000",53824 => "0000000000000000",
53825 => "0000000000000000",53826 => "0000000000000000",
53827 => "0000000000000000",53828 => "0000000000000000",
53829 => "0000000000000000",53830 => "0000000000000000",
53831 => "0000000000000000",53832 => "0000000000000000",
53833 => "0000000000000000",53834 => "0000000000000000",
53835 => "0000000000000000",53836 => "0000000000000000",
53837 => "0000000000000000",53838 => "0000000000000000",
53839 => "0000000000000000",53840 => "0000000000000000",
53841 => "0000000000000000",53842 => "0000000000000000",
53843 => "0000000000000000",53844 => "0000000000000000",
53845 => "0000000000000000",53846 => "0000000000000000",
53847 => "0000000000000000",53848 => "0000000000000000",
53849 => "0000000000000000",53850 => "0000000000000000",
53851 => "0000000000000000",53852 => "0000000000000000",
53853 => "0000000000000000",53854 => "0000000000000000",
53855 => "0000000000000000",53856 => "0000000000000000",
53857 => "0000000000000000",53858 => "0000000000000000",
53859 => "0000000000000000",53860 => "0000000000000000",
53861 => "0000000000000000",53862 => "0000000000000000",
53863 => "0000000000000000",53864 => "0000000000000000",
53865 => "0000000000000000",53866 => "0000000000000000",
53867 => "0000000000000000",53868 => "0000000000000000",
53869 => "0000000000000000",53870 => "0000000000000000",
53871 => "0000000000000000",53872 => "0000000000000000",
53873 => "0000000000000000",53874 => "0000000000000000",
53875 => "0000000000000000",53876 => "0000000000000000",
53877 => "0000000000000000",53878 => "0000000000000000",
53879 => "0000000000000000",53880 => "0000000000000000",
53881 => "0000000000000000",53882 => "0000000000000000",
53883 => "0000000000000000",53884 => "0000000000000000",
53885 => "0000000000000000",53886 => "0000000000000000",
53887 => "0000000000000000",53888 => "0000000000000000",
53889 => "0000000000000000",53890 => "0000000000000000",
53891 => "0000000000000000",53892 => "0000000000000000",
53893 => "0000000000000000",53894 => "0000000000000000",
53895 => "0000000000000000",53896 => "0000000000000000",
53897 => "0000000000000000",53898 => "0000000000000000",
53899 => "0000000000000000",53900 => "0000000000000000",
53901 => "0000000000000000",53902 => "0000000000000000",
53903 => "0000000000000000",53904 => "0000000000000000",
53905 => "0000000000000000",53906 => "0000000000000000",
53907 => "0000000000000000",53908 => "0000000000000000",
53909 => "0000000000000000",53910 => "0000000000000000",
53911 => "0000000000000000",53912 => "0000000000000000",
53913 => "0000000000000000",53914 => "0000000000000000",
53915 => "0000000000000000",53916 => "0000000000000000",
53917 => "0000000000000000",53918 => "0000000000000000",
53919 => "0000000000000000",53920 => "0000000000000000",
53921 => "0000000000000000",53922 => "0000000000000000",
53923 => "0000000000000000",53924 => "0000000000000000",
53925 => "0000000000000000",53926 => "0000000000000000",
53927 => "0000000000000000",53928 => "0000000000000000",
53929 => "0000000000000000",53930 => "0000000000000000",
53931 => "0000000000000000",53932 => "0000000000000000",
53933 => "0000000000000000",53934 => "0000000000000000",
53935 => "0000000000000000",53936 => "0000000000000000",
53937 => "0000000000000000",53938 => "0000000000000000",
53939 => "0000000000000000",53940 => "0000000000000000",
53941 => "0000000000000000",53942 => "0000000000000000",
53943 => "0000000000000000",53944 => "0000000000000000",
53945 => "0000000000000000",53946 => "0000000000000000",
53947 => "0000000000000000",53948 => "0000000000000000",
53949 => "0000000000000000",53950 => "0000000000000000",
53951 => "0000000000000000",53952 => "0000000000000000",
53953 => "0000000000000000",53954 => "0000000000000000",
53955 => "0000000000000000",53956 => "0000000000000000",
53957 => "0000000000000000",53958 => "0000000000000000",
53959 => "0000000000000000",53960 => "0000000000000000",
53961 => "0000000000000000",53962 => "0000000000000000",
53963 => "0000000000000000",53964 => "0000000000000000",
53965 => "0000000000000000",53966 => "0000000000000000",
53967 => "0000000000000000",53968 => "0000000000000000",
53969 => "0000000000000000",53970 => "0000000000000000",
53971 => "0000000000000000",53972 => "0000000000000000",
53973 => "0000000000000000",53974 => "0000000000000000",
53975 => "0000000000000000",53976 => "0000000000000000",
53977 => "0000000000000000",53978 => "0000000000000000",
53979 => "0000000000000000",53980 => "0000000000000000",
53981 => "0000000000000000",53982 => "0000000000000000",
53983 => "0000000000000000",53984 => "0000000000000000",
53985 => "0000000000000000",53986 => "0000000000000000",
53987 => "0000000000000000",53988 => "0000000000000000",
53989 => "0000000000000000",53990 => "0000000000000000",
53991 => "0000000000000000",53992 => "0000000000000000",
53993 => "0000000000000000",53994 => "0000000000000000",
53995 => "0000000000000000",53996 => "0000000000000000",
53997 => "0000000000000000",53998 => "0000000000000000",
53999 => "0000000000000000",54000 => "0000000000000000",
54001 => "0000000000000000",54002 => "0000000000000000",
54003 => "0000000000000000",54004 => "0000000000000000",
54005 => "0000000000000000",54006 => "0000000000000000",
54007 => "0000000000000000",54008 => "0000000000000000",
54009 => "0000000000000000",54010 => "0000000000000000",
54011 => "0000000000000000",54012 => "0000000000000000",
54013 => "0000000000000000",54014 => "0000000000000000",
54015 => "0000000000000000",54016 => "0000000000000000",
54017 => "0000000000000000",54018 => "0000000000000000",
54019 => "0000000000000000",54020 => "0000000000000000",
54021 => "0000000000000000",54022 => "0000000000000000",
54023 => "0000000000000000",54024 => "0000000000000000",
54025 => "0000000000000000",54026 => "0000000000000000",
54027 => "0000000000000000",54028 => "0000000000000000",
54029 => "0000000000000000",54030 => "0000000000000000",
54031 => "0000000000000000",54032 => "0000000000000000",
54033 => "0000000000000000",54034 => "0000000000000000",
54035 => "0000000000000000",54036 => "0000000000000000",
54037 => "0000000000000000",54038 => "0000000000000000",
54039 => "0000000000000000",54040 => "0000000000000000",
54041 => "0000000000000000",54042 => "0000000000000000",
54043 => "0000000000000000",54044 => "0000000000000000",
54045 => "0000000000000000",54046 => "0000000000000000",
54047 => "0000000000000000",54048 => "0000000000000000",
54049 => "0000000000000000",54050 => "0000000000000000",
54051 => "0000000000000000",54052 => "0000000000000000",
54053 => "0000000000000000",54054 => "0000000000000000",
54055 => "0000000000000000",54056 => "0000000000000000",
54057 => "0000000000000000",54058 => "0000000000000000",
54059 => "0000000000000000",54060 => "0000000000000000",
54061 => "0000000000000000",54062 => "0000000000000000",
54063 => "0000000000000000",54064 => "0000000000000000",
54065 => "0000000000000000",54066 => "0000000000000000",
54067 => "0000000000000000",54068 => "0000000000000000",
54069 => "0000000000000000",54070 => "0000000000000000",
54071 => "0000000000000000",54072 => "0000000000000000",
54073 => "0000000000000000",54074 => "0000000000000000",
54075 => "0000000000000000",54076 => "0000000000000000",
54077 => "0000000000000000",54078 => "0000000000000000",
54079 => "0000000000000000",54080 => "0000000000000000",
54081 => "0000000000000000",54082 => "0000000000000000",
54083 => "0000000000000000",54084 => "0000000000000000",
54085 => "0000000000000000",54086 => "0000000000000000",
54087 => "0000000000000000",54088 => "0000000000000000",
54089 => "0000000000000000",54090 => "0000000000000000",
54091 => "0000000000000000",54092 => "0000000000000000",
54093 => "0000000000000000",54094 => "0000000000000000",
54095 => "0000000000000000",54096 => "0000000000000000",
54097 => "0000000000000000",54098 => "0000000000000000",
54099 => "0000000000000000",54100 => "0000000000000000",
54101 => "0000000000000000",54102 => "0000000000000000",
54103 => "0000000000000000",54104 => "0000000000000000",
54105 => "0000000000000000",54106 => "0000000000000000",
54107 => "0000000000000000",54108 => "0000000000000000",
54109 => "0000000000000000",54110 => "0000000000000000",
54111 => "0000000000000000",54112 => "0000000000000000",
54113 => "0000000000000000",54114 => "0000000000000000",
54115 => "0000000000000000",54116 => "0000000000000000",
54117 => "0000000000000000",54118 => "0000000000000000",
54119 => "0000000000000000",54120 => "0000000000000000",
54121 => "0000000000000000",54122 => "0000000000000000",
54123 => "0000000000000000",54124 => "0000000000000000",
54125 => "0000000000000000",54126 => "0000000000000000",
54127 => "0000000000000000",54128 => "0000000000000000",
54129 => "0000000000000000",54130 => "0000000000000000",
54131 => "0000000000000000",54132 => "0000000000000000",
54133 => "0000000000000000",54134 => "0000000000000000",
54135 => "0000000000000000",54136 => "0000000000000000",
54137 => "0000000000000000",54138 => "0000000000000000",
54139 => "0000000000000000",54140 => "0000000000000000",
54141 => "0000000000000000",54142 => "0000000000000000",
54143 => "0000000000000000",54144 => "0000000000000000",
54145 => "0000000000000000",54146 => "0000000000000000",
54147 => "0000000000000000",54148 => "0000000000000000",
54149 => "0000000000000000",54150 => "0000000000000000",
54151 => "0000000000000000",54152 => "0000000000000000",
54153 => "0000000000000000",54154 => "0000000000000000",
54155 => "0000000000000000",54156 => "0000000000000000",
54157 => "0000000000000000",54158 => "0000000000000000",
54159 => "0000000000000000",54160 => "0000000000000000",
54161 => "0000000000000000",54162 => "0000000000000000",
54163 => "0000000000000000",54164 => "0000000000000000",
54165 => "0000000000000000",54166 => "0000000000000000",
54167 => "0000000000000000",54168 => "0000000000000000",
54169 => "0000000000000000",54170 => "0000000000000000",
54171 => "0000000000000000",54172 => "0000000000000000",
54173 => "0000000000000000",54174 => "0000000000000000",
54175 => "0000000000000000",54176 => "0000000000000000",
54177 => "0000000000000000",54178 => "0000000000000000",
54179 => "0000000000000000",54180 => "0000000000000000",
54181 => "0000000000000000",54182 => "0000000000000000",
54183 => "0000000000000000",54184 => "0000000000000000",
54185 => "0000000000000000",54186 => "0000000000000000",
54187 => "0000000000000000",54188 => "0000000000000000",
54189 => "0000000000000000",54190 => "0000000000000000",
54191 => "0000000000000000",54192 => "0000000000000000",
54193 => "0000000000000000",54194 => "0000000000000000",
54195 => "0000000000000000",54196 => "0000000000000000",
54197 => "0000000000000000",54198 => "0000000000000000",
54199 => "0000000000000000",54200 => "0000000000000000",
54201 => "0000000000000000",54202 => "0000000000000000",
54203 => "0000000000000000",54204 => "0000000000000000",
54205 => "0000000000000000",54206 => "0000000000000000",
54207 => "0000000000000000",54208 => "0000000000000000",
54209 => "0000000000000000",54210 => "0000000000000000",
54211 => "0000000000000000",54212 => "0000000000000000",
54213 => "0000000000000000",54214 => "0000000000000000",
54215 => "0000000000000000",54216 => "0000000000000000",
54217 => "0000000000000000",54218 => "0000000000000000",
54219 => "0000000000000000",54220 => "0000000000000000",
54221 => "0000000000000000",54222 => "0000000000000000",
54223 => "0000000000000000",54224 => "0000000000000000",
54225 => "0000000000000000",54226 => "0000000000000000",
54227 => "0000000000000000",54228 => "0000000000000000",
54229 => "0000000000000000",54230 => "0000000000000000",
54231 => "0000000000000000",54232 => "0000000000000000",
54233 => "0000000000000000",54234 => "0000000000000000",
54235 => "0000000000000000",54236 => "0000000000000000",
54237 => "0000000000000000",54238 => "0000000000000000",
54239 => "0000000000000000",54240 => "0000000000000000",
54241 => "0000000000000000",54242 => "0000000000000000",
54243 => "0000000000000000",54244 => "0000000000000000",
54245 => "0000000000000000",54246 => "0000000000000000",
54247 => "0000000000000000",54248 => "0000000000000000",
54249 => "0000000000000000",54250 => "0000000000000000",
54251 => "0000000000000000",54252 => "0000000000000000",
54253 => "0000000000000000",54254 => "0000000000000000",
54255 => "0000000000000000",54256 => "0000000000000000",
54257 => "0000000000000000",54258 => "0000000000000000",
54259 => "0000000000000000",54260 => "0000000000000000",
54261 => "0000000000000000",54262 => "0000000000000000",
54263 => "0000000000000000",54264 => "0000000000000000",
54265 => "0000000000000000",54266 => "0000000000000000",
54267 => "0000000000000000",54268 => "0000000000000000",
54269 => "0000000000000000",54270 => "0000000000000000",
54271 => "0000000000000000",54272 => "0000000000000000",
54273 => "0000000000000000",54274 => "0000000000000000",
54275 => "0000000000000000",54276 => "0000000000000000",
54277 => "0000000000000000",54278 => "0000000000000000",
54279 => "0000000000000000",54280 => "0000000000000000",
54281 => "0000000000000000",54282 => "0000000000000000",
54283 => "0000000000000000",54284 => "0000000000000000",
54285 => "0000000000000000",54286 => "0000000000000000",
54287 => "0000000000000000",54288 => "0000000000000000",
54289 => "0000000000000000",54290 => "0000000000000000",
54291 => "0000000000000000",54292 => "0000000000000000",
54293 => "0000000000000000",54294 => "0000000000000000",
54295 => "0000000000000000",54296 => "0000000000000000",
54297 => "0000000000000000",54298 => "0000000000000000",
54299 => "0000000000000000",54300 => "0000000000000000",
54301 => "0000000000000000",54302 => "0000000000000000",
54303 => "0000000000000000",54304 => "0000000000000000",
54305 => "0000000000000000",54306 => "0000000000000000",
54307 => "0000000000000000",54308 => "0000000000000000",
54309 => "0000000000000000",54310 => "0000000000000000",
54311 => "0000000000000000",54312 => "0000000000000000",
54313 => "0000000000000000",54314 => "0000000000000000",
54315 => "0000000000000000",54316 => "0000000000000000",
54317 => "0000000000000000",54318 => "0000000000000000",
54319 => "0000000000000000",54320 => "0000000000000000",
54321 => "0000000000000000",54322 => "0000000000000000",
54323 => "0000000000000000",54324 => "0000000000000000",
54325 => "0000000000000000",54326 => "0000000000000000",
54327 => "0000000000000000",54328 => "0000000000000000",
54329 => "0000000000000000",54330 => "0000000000000000",
54331 => "0000000000000000",54332 => "0000000000000000",
54333 => "0000000000000000",54334 => "0000000000000000",
54335 => "0000000000000000",54336 => "0000000000000000",
54337 => "0000000000000000",54338 => "0000000000000000",
54339 => "0000000000000000",54340 => "0000000000000000",
54341 => "0000000000000000",54342 => "0000000000000000",
54343 => "0000000000000000",54344 => "0000000000000000",
54345 => "0000000000000000",54346 => "0000000000000000",
54347 => "0000000000000000",54348 => "0000000000000000",
54349 => "0000000000000000",54350 => "0000000000000000",
54351 => "0000000000000000",54352 => "0000000000000000",
54353 => "0000000000000000",54354 => "0000000000000000",
54355 => "0000000000000000",54356 => "0000000000000000",
54357 => "0000000000000000",54358 => "0000000000000000",
54359 => "0000000000000000",54360 => "0000000000000000",
54361 => "0000000000000000",54362 => "0000000000000000",
54363 => "0000000000000000",54364 => "0000000000000000",
54365 => "0000000000000000",54366 => "0000000000000000",
54367 => "0000000000000000",54368 => "0000000000000000",
54369 => "0000000000000000",54370 => "0000000000000000",
54371 => "0000000000000000",54372 => "0000000000000000",
54373 => "0000000000000000",54374 => "0000000000000000",
54375 => "0000000000000000",54376 => "0000000000000000",
54377 => "0000000000000000",54378 => "0000000000000000",
54379 => "0000000000000000",54380 => "0000000000000000",
54381 => "0000000000000000",54382 => "0000000000000000",
54383 => "0000000000000000",54384 => "0000000000000000",
54385 => "0000000000000000",54386 => "0000000000000000",
54387 => "0000000000000000",54388 => "0000000000000000",
54389 => "0000000000000000",54390 => "0000000000000000",
54391 => "0000000000000000",54392 => "0000000000000000",
54393 => "0000000000000000",54394 => "0000000000000000",
54395 => "0000000000000000",54396 => "0000000000000000",
54397 => "0000000000000000",54398 => "0000000000000000",
54399 => "0000000000000000",54400 => "0000000000000000",
54401 => "0000000000000000",54402 => "0000000000000000",
54403 => "0000000000000000",54404 => "0000000000000000",
54405 => "0000000000000000",54406 => "0000000000000000",
54407 => "0000000000000000",54408 => "0000000000000000",
54409 => "0000000000000000",54410 => "0000000000000000",
54411 => "0000000000000000",54412 => "0000000000000000",
54413 => "0000000000000000",54414 => "0000000000000000",
54415 => "0000000000000000",54416 => "0000000000000000",
54417 => "0000000000000000",54418 => "0000000000000000",
54419 => "0000000000000000",54420 => "0000000000000000",
54421 => "0000000000000000",54422 => "0000000000000000",
54423 => "0000000000000000",54424 => "0000000000000000",
54425 => "0000000000000000",54426 => "0000000000000000",
54427 => "0000000000000000",54428 => "0000000000000000",
54429 => "0000000000000000",54430 => "0000000000000000",
54431 => "0000000000000000",54432 => "0000000000000000",
54433 => "0000000000000000",54434 => "0000000000000000",
54435 => "0000000000000000",54436 => "0000000000000000",
54437 => "0000000000000000",54438 => "0000000000000000",
54439 => "0000000000000000",54440 => "0000000000000000",
54441 => "0000000000000000",54442 => "0000000000000000",
54443 => "0000000000000000",54444 => "0000000000000000",
54445 => "0000000000000000",54446 => "0000000000000000",
54447 => "0000000000000000",54448 => "0000000000000000",
54449 => "0000000000000000",54450 => "0000000000000000",
54451 => "0000000000000000",54452 => "0000000000000000",
54453 => "0000000000000000",54454 => "0000000000000000",
54455 => "0000000000000000",54456 => "0000000000000000",
54457 => "0000000000000000",54458 => "0000000000000000",
54459 => "0000000000000000",54460 => "0000000000000000",
54461 => "0000000000000000",54462 => "0000000000000000",
54463 => "0000000000000000",54464 => "0000000000000000",
54465 => "0000000000000000",54466 => "0000000000000000",
54467 => "0000000000000000",54468 => "0000000000000000",
54469 => "0000000000000000",54470 => "0000000000000000",
54471 => "0000000000000000",54472 => "0000000000000000",
54473 => "0000000000000000",54474 => "0000000000000000",
54475 => "0000000000000000",54476 => "0000000000000000",
54477 => "0000000000000000",54478 => "0000000000000000",
54479 => "0000000000000000",54480 => "0000000000000000",
54481 => "0000000000000000",54482 => "0000000000000000",
54483 => "0000000000000000",54484 => "0000000000000000",
54485 => "0000000000000000",54486 => "0000000000000000",
54487 => "0000000000000000",54488 => "0000000000000000",
54489 => "0000000000000000",54490 => "0000000000000000",
54491 => "0000000000000000",54492 => "0000000000000000",
54493 => "0000000000000000",54494 => "0000000000000000",
54495 => "0000000000000000",54496 => "0000000000000000",
54497 => "0000000000000000",54498 => "0000000000000000",
54499 => "0000000000000000",54500 => "0000000000000000",
54501 => "0000000000000000",54502 => "0000000000000000",
54503 => "0000000000000000",54504 => "0000000000000000",
54505 => "0000000000000000",54506 => "0000000000000000",
54507 => "0000000000000000",54508 => "0000000000000000",
54509 => "0000000000000000",54510 => "0000000000000000",
54511 => "0000000000000000",54512 => "0000000000000000",
54513 => "0000000000000000",54514 => "0000000000000000",
54515 => "0000000000000000",54516 => "0000000000000000",
54517 => "0000000000000000",54518 => "0000000000000000",
54519 => "0000000000000000",54520 => "0000000000000000",
54521 => "0000000000000000",54522 => "0000000000000000",
54523 => "0000000000000000",54524 => "0000000000000000",
54525 => "0000000000000000",54526 => "0000000000000000",
54527 => "0000000000000000",54528 => "0000000000000000",
54529 => "0000000000000000",54530 => "0000000000000000",
54531 => "0000000000000000",54532 => "0000000000000000",
54533 => "0000000000000000",54534 => "0000000000000000",
54535 => "0000000000000000",54536 => "0000000000000000",
54537 => "0000000000000000",54538 => "0000000000000000",
54539 => "0000000000000000",54540 => "0000000000000000",
54541 => "0000000000000000",54542 => "0000000000000000",
54543 => "0000000000000000",54544 => "0000000000000000",
54545 => "0000000000000000",54546 => "0000000000000000",
54547 => "0000000000000000",54548 => "0000000000000000",
54549 => "0000000000000000",54550 => "0000000000000000",
54551 => "0000000000000000",54552 => "0000000000000000",
54553 => "0000000000000000",54554 => "0000000000000000",
54555 => "0000000000000000",54556 => "0000000000000000",
54557 => "0000000000000000",54558 => "0000000000000000",
54559 => "0000000000000000",54560 => "0000000000000000",
54561 => "0000000000000000",54562 => "0000000000000000",
54563 => "0000000000000000",54564 => "0000000000000000",
54565 => "0000000000000000",54566 => "0000000000000000",
54567 => "0000000000000000",54568 => "0000000000000000",
54569 => "0000000000000000",54570 => "0000000000000000",
54571 => "0000000000000000",54572 => "0000000000000000",
54573 => "0000000000000000",54574 => "0000000000000000",
54575 => "0000000000000000",54576 => "0000000000000000",
54577 => "0000000000000000",54578 => "0000000000000000",
54579 => "0000000000000000",54580 => "0000000000000000",
54581 => "0000000000000000",54582 => "0000000000000000",
54583 => "0000000000000000",54584 => "0000000000000000",
54585 => "0000000000000000",54586 => "0000000000000000",
54587 => "0000000000000000",54588 => "0000000000000000",
54589 => "0000000000000000",54590 => "0000000000000000",
54591 => "0000000000000000",54592 => "0000000000000000",
54593 => "0000000000000000",54594 => "0000000000000000",
54595 => "0000000000000000",54596 => "0000000000000000",
54597 => "0000000000000000",54598 => "0000000000000000",
54599 => "0000000000000000",54600 => "0000000000000000",
54601 => "0000000000000000",54602 => "0000000000000000",
54603 => "0000000000000000",54604 => "0000000000000000",
54605 => "0000000000000000",54606 => "0000000000000000",
54607 => "0000000000000000",54608 => "0000000000000000",
54609 => "0000000000000000",54610 => "0000000000000000",
54611 => "0000000000000000",54612 => "0000000000000000",
54613 => "0000000000000000",54614 => "0000000000000000",
54615 => "0000000000000000",54616 => "0000000000000000",
54617 => "0000000000000000",54618 => "0000000000000000",
54619 => "0000000000000000",54620 => "0000000000000000",
54621 => "0000000000000000",54622 => "0000000000000000",
54623 => "0000000000000000",54624 => "0000000000000000",
54625 => "0000000000000000",54626 => "0000000000000000",
54627 => "0000000000000000",54628 => "0000000000000000",
54629 => "0000000000000000",54630 => "0000000000000000",
54631 => "0000000000000000",54632 => "0000000000000000",
54633 => "0000000000000000",54634 => "0000000000000000",
54635 => "0000000000000000",54636 => "0000000000000000",
54637 => "0000000000000000",54638 => "0000000000000000",
54639 => "0000000000000000",54640 => "0000000000000000",
54641 => "0000000000000000",54642 => "0000000000000000",
54643 => "0000000000000000",54644 => "0000000000000000",
54645 => "0000000000000000",54646 => "0000000000000000",
54647 => "0000000000000000",54648 => "0000000000000000",
54649 => "0000000000000000",54650 => "0000000000000000",
54651 => "0000000000000000",54652 => "0000000000000000",
54653 => "0000000000000000",54654 => "0000000000000000",
54655 => "0000000000000000",54656 => "0000000000000000",
54657 => "0000000000000000",54658 => "0000000000000000",
54659 => "0000000000000000",54660 => "0000000000000000",
54661 => "0000000000000000",54662 => "0000000000000000",
54663 => "0000000000000000",54664 => "0000000000000000",
54665 => "0000000000000000",54666 => "0000000000000000",
54667 => "0000000000000000",54668 => "0000000000000000",
54669 => "0000000000000000",54670 => "0000000000000000",
54671 => "0000000000000000",54672 => "0000000000000000",
54673 => "0000000000000000",54674 => "0000000000000000",
54675 => "0000000000000000",54676 => "0000000000000000",
54677 => "0000000000000000",54678 => "0000000000000000",
54679 => "0000000000000000",54680 => "0000000000000000",
54681 => "0000000000000000",54682 => "0000000000000000",
54683 => "0000000000000000",54684 => "0000000000000000",
54685 => "0000000000000000",54686 => "0000000000000000",
54687 => "0000000000000000",54688 => "0000000000000000",
54689 => "0000000000000000",54690 => "0000000000000000",
54691 => "0000000000000000",54692 => "0000000000000000",
54693 => "0000000000000000",54694 => "0000000000000000",
54695 => "0000000000000000",54696 => "0000000000000000",
54697 => "0000000000000000",54698 => "0000000000000000",
54699 => "0000000000000000",54700 => "0000000000000000",
54701 => "0000000000000000",54702 => "0000000000000000",
54703 => "0000000000000000",54704 => "0000000000000000",
54705 => "0000000000000000",54706 => "0000000000000000",
54707 => "0000000000000000",54708 => "0000000000000000",
54709 => "0000000000000000",54710 => "0000000000000000",
54711 => "0000000000000000",54712 => "0000000000000000",
54713 => "0000000000000000",54714 => "0000000000000000",
54715 => "0000000000000000",54716 => "0000000000000000",
54717 => "0000000000000000",54718 => "0000000000000000",
54719 => "0000000000000000",54720 => "0000000000000000",
54721 => "0000000000000000",54722 => "0000000000000000",
54723 => "0000000000000000",54724 => "0000000000000000",
54725 => "0000000000000000",54726 => "0000000000000000",
54727 => "0000000000000000",54728 => "0000000000000000",
54729 => "0000000000000000",54730 => "0000000000000000",
54731 => "0000000000000000",54732 => "0000000000000000",
54733 => "0000000000000000",54734 => "0000000000000000",
54735 => "0000000000000000",54736 => "0000000000000000",
54737 => "0000000000000000",54738 => "0000000000000000",
54739 => "0000000000000000",54740 => "0000000000000000",
54741 => "0000000000000000",54742 => "0000000000000000",
54743 => "0000000000000000",54744 => "0000000000000000",
54745 => "0000000000000000",54746 => "0000000000000000",
54747 => "0000000000000000",54748 => "0000000000000000",
54749 => "0000000000000000",54750 => "0000000000000000",
54751 => "0000000000000000",54752 => "0000000000000000",
54753 => "0000000000000000",54754 => "0000000000000000",
54755 => "0000000000000000",54756 => "0000000000000000",
54757 => "0000000000000000",54758 => "0000000000000000",
54759 => "0000000000000000",54760 => "0000000000000000",
54761 => "0000000000000000",54762 => "0000000000000000",
54763 => "0000000000000000",54764 => "0000000000000000",
54765 => "0000000000000000",54766 => "0000000000000000",
54767 => "0000000000000000",54768 => "0000000000000000",
54769 => "0000000000000000",54770 => "0000000000000000",
54771 => "0000000000000000",54772 => "0000000000000000",
54773 => "0000000000000000",54774 => "0000000000000000",
54775 => "0000000000000000",54776 => "0000000000000000",
54777 => "0000000000000000",54778 => "0000000000000000",
54779 => "0000000000000000",54780 => "0000000000000000",
54781 => "0000000000000000",54782 => "0000000000000000",
54783 => "0000000000000000",54784 => "0000000000000000",
54785 => "0000000000000000",54786 => "0000000000000000",
54787 => "0000000000000000",54788 => "0000000000000000",
54789 => "0000000000000000",54790 => "0000000000000000",
54791 => "0000000000000000",54792 => "0000000000000000",
54793 => "0000000000000000",54794 => "0000000000000000",
54795 => "0000000000000000",54796 => "0000000000000000",
54797 => "0000000000000000",54798 => "0000000000000000",
54799 => "0000000000000000",54800 => "0000000000000000",
54801 => "0000000000000000",54802 => "0000000000000000",
54803 => "0000000000000000",54804 => "0000000000000000",
54805 => "0000000000000000",54806 => "0000000000000000",
54807 => "0000000000000000",54808 => "0000000000000000",
54809 => "0000000000000000",54810 => "0000000000000000",
54811 => "0000000000000000",54812 => "0000000000000000",
54813 => "0000000000000000",54814 => "0000000000000000",
54815 => "0000000000000000",54816 => "0000000000000000",
54817 => "0000000000000000",54818 => "0000000000000000",
54819 => "0000000000000000",54820 => "0000000000000000",
54821 => "0000000000000000",54822 => "0000000000000000",
54823 => "0000000000000000",54824 => "0000000000000000",
54825 => "0000000000000000",54826 => "0000000000000000",
54827 => "0000000000000000",54828 => "0000000000000000",
54829 => "0000000000000000",54830 => "0000000000000000",
54831 => "0000000000000000",54832 => "0000000000000000",
54833 => "0000000000000000",54834 => "0000000000000000",
54835 => "0000000000000000",54836 => "0000000000000000",
54837 => "0000000000000000",54838 => "0000000000000000",
54839 => "0000000000000000",54840 => "0000000000000000",
54841 => "0000000000000000",54842 => "0000000000000000",
54843 => "0000000000000000",54844 => "0000000000000000",
54845 => "0000000000000000",54846 => "0000000000000000",
54847 => "0000000000000000",54848 => "0000000000000000",
54849 => "0000000000000000",54850 => "0000000000000000",
54851 => "0000000000000000",54852 => "0000000000000000",
54853 => "0000000000000000",54854 => "0000000000000000",
54855 => "0000000000000000",54856 => "0000000000000000",
54857 => "0000000000000000",54858 => "0000000000000000",
54859 => "0000000000000000",54860 => "0000000000000000",
54861 => "0000000000000000",54862 => "0000000000000000",
54863 => "0000000000000000",54864 => "0000000000000000",
54865 => "0000000000000000",54866 => "0000000000000000",
54867 => "0000000000000000",54868 => "0000000000000000",
54869 => "0000000000000000",54870 => "0000000000000000",
54871 => "0000000000000000",54872 => "0000000000000000",
54873 => "0000000000000000",54874 => "0000000000000000",
54875 => "0000000000000000",54876 => "0000000000000000",
54877 => "0000000000000000",54878 => "0000000000000000",
54879 => "0000000000000000",54880 => "0000000000000000",
54881 => "0000000000000000",54882 => "0000000000000000",
54883 => "0000000000000000",54884 => "0000000000000000",
54885 => "0000000000000000",54886 => "0000000000000000",
54887 => "0000000000000000",54888 => "0000000000000000",
54889 => "0000000000000000",54890 => "0000000000000000",
54891 => "0000000000000000",54892 => "0000000000000000",
54893 => "0000000000000000",54894 => "0000000000000000",
54895 => "0000000000000000",54896 => "0000000000000000",
54897 => "0000000000000000",54898 => "0000000000000000",
54899 => "0000000000000000",54900 => "0000000000000000",
54901 => "0000000000000000",54902 => "0000000000000000",
54903 => "0000000000000000",54904 => "0000000000000000",
54905 => "0000000000000000",54906 => "0000000000000000",
54907 => "0000000000000000",54908 => "0000000000000000",
54909 => "0000000000000000",54910 => "0000000000000000",
54911 => "0000000000000000",54912 => "0000000000000000",
54913 => "0000000000000000",54914 => "0000000000000000",
54915 => "0000000000000000",54916 => "0000000000000000",
54917 => "0000000000000000",54918 => "0000000000000000",
54919 => "0000000000000000",54920 => "0000000000000000",
54921 => "0000000000000000",54922 => "0000000000000000",
54923 => "0000000000000000",54924 => "0000000000000000",
54925 => "0000000000000000",54926 => "0000000000000000",
54927 => "0000000000000000",54928 => "0000000000000000",
54929 => "0000000000000000",54930 => "0000000000000000",
54931 => "0000000000000000",54932 => "0000000000000000",
54933 => "0000000000000000",54934 => "0000000000000000",
54935 => "0000000000000000",54936 => "0000000000000000",
54937 => "0000000000000000",54938 => "0000000000000000",
54939 => "0000000000000000",54940 => "0000000000000000",
54941 => "0000000000000000",54942 => "0000000000000000",
54943 => "0000000000000000",54944 => "0000000000000000",
54945 => "0000000000000000",54946 => "0000000000000000",
54947 => "0000000000000000",54948 => "0000000000000000",
54949 => "0000000000000000",54950 => "0000000000000000",
54951 => "0000000000000000",54952 => "0000000000000000",
54953 => "0000000000000000",54954 => "0000000000000000",
54955 => "0000000000000000",54956 => "0000000000000000",
54957 => "0000000000000000",54958 => "0000000000000000",
54959 => "0000000000000000",54960 => "0000000000000000",
54961 => "0000000000000000",54962 => "0000000000000000",
54963 => "0000000000000000",54964 => "0000000000000000",
54965 => "0000000000000000",54966 => "0000000000000000",
54967 => "0000000000000000",54968 => "0000000000000000",
54969 => "0000000000000000",54970 => "0000000000000000",
54971 => "0000000000000000",54972 => "0000000000000000",
54973 => "0000000000000000",54974 => "0000000000000000",
54975 => "0000000000000000",54976 => "0000000000000000",
54977 => "0000000000000000",54978 => "0000000000000000",
54979 => "0000000000000000",54980 => "0000000000000000",
54981 => "0000000000000000",54982 => "0000000000000000",
54983 => "0000000000000000",54984 => "0000000000000000",
54985 => "0000000000000000",54986 => "0000000000000000",
54987 => "0000000000000000",54988 => "0000000000000000",
54989 => "0000000000000000",54990 => "0000000000000000",
54991 => "0000000000000000",54992 => "0000000000000000",
54993 => "0000000000000000",54994 => "0000000000000000",
54995 => "0000000000000000",54996 => "0000000000000000",
54997 => "0000000000000000",54998 => "0000000000000000",
54999 => "0000000000000000",55000 => "0000000000000000",
55001 => "0000000000000000",55002 => "0000000000000000",
55003 => "0000000000000000",55004 => "0000000000000000",
55005 => "0000000000000000",55006 => "0000000000000000",
55007 => "0000000000000000",55008 => "0000000000000000",
55009 => "0000000000000000",55010 => "0000000000000000",
55011 => "0000000000000000",55012 => "0000000000000000",
55013 => "0000000000000000",55014 => "0000000000000000",
55015 => "0000000000000000",55016 => "0000000000000000",
55017 => "0000000000000000",55018 => "0000000000000000",
55019 => "0000000000000000",55020 => "0000000000000000",
55021 => "0000000000000000",55022 => "0000000000000000",
55023 => "0000000000000000",55024 => "0000000000000000",
55025 => "0000000000000000",55026 => "0000000000000000",
55027 => "0000000000000000",55028 => "0000000000000000",
55029 => "0000000000000000",55030 => "0000000000000000",
55031 => "0000000000000000",55032 => "0000000000000000",
55033 => "0000000000000000",55034 => "0000000000000000",
55035 => "0000000000000000",55036 => "0000000000000000",
55037 => "0000000000000000",55038 => "0000000000000000",
55039 => "0000000000000000",55040 => "0000000000000000",
55041 => "0000000000000000",55042 => "0000000000000000",
55043 => "0000000000000000",55044 => "0000000000000000",
55045 => "0000000000000000",55046 => "0000000000000000",
55047 => "0000000000000000",55048 => "0000000000000000",
55049 => "0000000000000000",55050 => "0000000000000000",
55051 => "0000000000000000",55052 => "0000000000000000",
55053 => "0000000000000000",55054 => "0000000000000000",
55055 => "0000000000000000",55056 => "0000000000000000",
55057 => "0000000000000000",55058 => "0000000000000000",
55059 => "0000000000000000",55060 => "0000000000000000",
55061 => "0000000000000000",55062 => "0000000000000000",
55063 => "0000000000000000",55064 => "0000000000000000",
55065 => "0000000000000000",55066 => "0000000000000000",
55067 => "0000000000000000",55068 => "0000000000000000",
55069 => "0000000000000000",55070 => "0000000000000000",
55071 => "0000000000000000",55072 => "0000000000000000",
55073 => "0000000000000000",55074 => "0000000000000000",
55075 => "0000000000000000",55076 => "0000000000000000",
55077 => "0000000000000000",55078 => "0000000000000000",
55079 => "0000000000000000",55080 => "0000000000000000",
55081 => "0000000000000000",55082 => "0000000000000000",
55083 => "0000000000000000",55084 => "0000000000000000",
55085 => "0000000000000000",55086 => "0000000000000000",
55087 => "0000000000000000",55088 => "0000000000000000",
55089 => "0000000000000000",55090 => "0000000000000000",
55091 => "0000000000000000",55092 => "0000000000000000",
55093 => "0000000000000000",55094 => "0000000000000000",
55095 => "0000000000000000",55096 => "0000000000000000",
55097 => "0000000000000000",55098 => "0000000000000000",
55099 => "0000000000000000",55100 => "0000000000000000",
55101 => "0000000000000000",55102 => "0000000000000000",
55103 => "0000000000000000",55104 => "0000000000000000",
55105 => "0000000000000000",55106 => "0000000000000000",
55107 => "0000000000000000",55108 => "0000000000000000",
55109 => "0000000000000000",55110 => "0000000000000000",
55111 => "0000000000000000",55112 => "0000000000000000",
55113 => "0000000000000000",55114 => "0000000000000000",
55115 => "0000000000000000",55116 => "0000000000000000",
55117 => "0000000000000000",55118 => "0000000000000000",
55119 => "0000000000000000",55120 => "0000000000000000",
55121 => "0000000000000000",55122 => "0000000000000000",
55123 => "0000000000000000",55124 => "0000000000000000",
55125 => "0000000000000000",55126 => "0000000000000000",
55127 => "0000000000000000",55128 => "0000000000000000",
55129 => "0000000000000000",55130 => "0000000000000000",
55131 => "0000000000000000",55132 => "0000000000000000",
55133 => "0000000000000000",55134 => "0000000000000000",
55135 => "0000000000000000",55136 => "0000000000000000",
55137 => "0000000000000000",55138 => "0000000000000000",
55139 => "0000000000000000",55140 => "0000000000000000",
55141 => "0000000000000000",55142 => "0000000000000000",
55143 => "0000000000000000",55144 => "0000000000000000",
55145 => "0000000000000000",55146 => "0000000000000000",
55147 => "0000000000000000",55148 => "0000000000000000",
55149 => "0000000000000000",55150 => "0000000000000000",
55151 => "0000000000000000",55152 => "0000000000000000",
55153 => "0000000000000000",55154 => "0000000000000000",
55155 => "0000000000000000",55156 => "0000000000000000",
55157 => "0000000000000000",55158 => "0000000000000000",
55159 => "0000000000000000",55160 => "0000000000000000",
55161 => "0000000000000000",55162 => "0000000000000000",
55163 => "0000000000000000",55164 => "0000000000000000",
55165 => "0000000000000000",55166 => "0000000000000000",
55167 => "0000000000000000",55168 => "0000000000000000",
55169 => "0000000000000000",55170 => "0000000000000000",
55171 => "0000000000000000",55172 => "0000000000000000",
55173 => "0000000000000000",55174 => "0000000000000000",
55175 => "0000000000000000",55176 => "0000000000000000",
55177 => "0000000000000000",55178 => "0000000000000000",
55179 => "0000000000000000",55180 => "0000000000000000",
55181 => "0000000000000000",55182 => "0000000000000000",
55183 => "0000000000000000",55184 => "0000000000000000",
55185 => "0000000000000000",55186 => "0000000000000000",
55187 => "0000000000000000",55188 => "0000000000000000",
55189 => "0000000000000000",55190 => "0000000000000000",
55191 => "0000000000000000",55192 => "0000000000000000",
55193 => "0000000000000000",55194 => "0000000000000000",
55195 => "0000000000000000",55196 => "0000000000000000",
55197 => "0000000000000000",55198 => "0000000000000000",
55199 => "0000000000000000",55200 => "0000000000000000",
55201 => "0000000000000000",55202 => "0000000000000000",
55203 => "0000000000000000",55204 => "0000000000000000",
55205 => "0000000000000000",55206 => "0000000000000000",
55207 => "0000000000000000",55208 => "0000000000000000",
55209 => "0000000000000000",55210 => "0000000000000000",
55211 => "0000000000000000",55212 => "0000000000000000",
55213 => "0000000000000000",55214 => "0000000000000000",
55215 => "0000000000000000",55216 => "0000000000000000",
55217 => "0000000000000000",55218 => "0000000000000000",
55219 => "0000000000000000",55220 => "0000000000000000",
55221 => "0000000000000000",55222 => "0000000000000000",
55223 => "0000000000000000",55224 => "0000000000000000",
55225 => "0000000000000000",55226 => "0000000000000000",
55227 => "0000000000000000",55228 => "0000000000000000",
55229 => "0000000000000000",55230 => "0000000000000000",
55231 => "0000000000000000",55232 => "0000000000000000",
55233 => "0000000000000000",55234 => "0000000000000000",
55235 => "0000000000000000",55236 => "0000000000000000",
55237 => "0000000000000000",55238 => "0000000000000000",
55239 => "0000000000000000",55240 => "0000000000000000",
55241 => "0000000000000000",55242 => "0000000000000000",
55243 => "0000000000000000",55244 => "0000000000000000",
55245 => "0000000000000000",55246 => "0000000000000000",
55247 => "0000000000000000",55248 => "0000000000000000",
55249 => "0000000000000000",55250 => "0000000000000000",
55251 => "0000000000000000",55252 => "0000000000000000",
55253 => "0000000000000000",55254 => "0000000000000000",
55255 => "0000000000000000",55256 => "0000000000000000",
55257 => "0000000000000000",55258 => "0000000000000000",
55259 => "0000000000000000",55260 => "0000000000000000",
55261 => "0000000000000000",55262 => "0000000000000000",
55263 => "0000000000000000",55264 => "0000000000000000",
55265 => "0000000000000000",55266 => "0000000000000000",
55267 => "0000000000000000",55268 => "0000000000000000",
55269 => "0000000000000000",55270 => "0000000000000000",
55271 => "0000000000000000",55272 => "0000000000000000",
55273 => "0000000000000000",55274 => "0000000000000000",
55275 => "0000000000000000",55276 => "0000000000000000",
55277 => "0000000000000000",55278 => "0000000000000000",
55279 => "0000000000000000",55280 => "0000000000000000",
55281 => "0000000000000000",55282 => "0000000000000000",
55283 => "0000000000000000",55284 => "0000000000000000",
55285 => "0000000000000000",55286 => "0000000000000000",
55287 => "0000000000000000",55288 => "0000000000000000",
55289 => "0000000000000000",55290 => "0000000000000000",
55291 => "0000000000000000",55292 => "0000000000000000",
55293 => "0000000000000000",55294 => "0000000000000000",
55295 => "0000000000000000",55296 => "0000000000000000",
55297 => "0000000000000000",55298 => "0000000000000000",
55299 => "0000000000000000",55300 => "0000000000000000",
55301 => "0000000000000000",55302 => "0000000000000000",
55303 => "0000000000000000",55304 => "0000000000000000",
55305 => "0000000000000000",55306 => "0000000000000000",
55307 => "0000000000000000",55308 => "0000000000000000",
55309 => "0000000000000000",55310 => "0000000000000000",
55311 => "0000000000000000",55312 => "0000000000000000",
55313 => "0000000000000000",55314 => "0000000000000000",
55315 => "0000000000000000",55316 => "0000000000000000",
55317 => "0000000000000000",55318 => "0000000000000000",
55319 => "0000000000000000",55320 => "0000000000000000",
55321 => "0000000000000000",55322 => "0000000000000000",
55323 => "0000000000000000",55324 => "0000000000000000",
55325 => "0000000000000000",55326 => "0000000000000000",
55327 => "0000000000000000",55328 => "0000000000000000",
55329 => "0000000000000000",55330 => "0000000000000000",
55331 => "0000000000000000",55332 => "0000000000000000",
55333 => "0000000000000000",55334 => "0000000000000000",
55335 => "0000000000000000",55336 => "0000000000000000",
55337 => "0000000000000000",55338 => "0000000000000000",
55339 => "0000000000000000",55340 => "0000000000000000",
55341 => "0000000000000000",55342 => "0000000000000000",
55343 => "0000000000000000",55344 => "0000000000000000",
55345 => "0000000000000000",55346 => "0000000000000000",
55347 => "0000000000000000",55348 => "0000000000000000",
55349 => "0000000000000000",55350 => "0000000000000000",
55351 => "0000000000000000",55352 => "0000000000000000",
55353 => "0000000000000000",55354 => "0000000000000000",
55355 => "0000000000000000",55356 => "0000000000000000",
55357 => "0000000000000000",55358 => "0000000000000000",
55359 => "0000000000000000",55360 => "0000000000000000",
55361 => "0000000000000000",55362 => "0000000000000000",
55363 => "0000000000000000",55364 => "0000000000000000",
55365 => "0000000000000000",55366 => "0000000000000000",
55367 => "0000000000000000",55368 => "0000000000000000",
55369 => "0000000000000000",55370 => "0000000000000000",
55371 => "0000000000000000",55372 => "0000000000000000",
55373 => "0000000000000000",55374 => "0000000000000000",
55375 => "0000000000000000",55376 => "0000000000000000",
55377 => "0000000000000000",55378 => "0000000000000000",
55379 => "0000000000000000",55380 => "0000000000000000",
55381 => "0000000000000000",55382 => "0000000000000000",
55383 => "0000000000000000",55384 => "0000000000000000",
55385 => "0000000000000000",55386 => "0000000000000000",
55387 => "0000000000000000",55388 => "0000000000000000",
55389 => "0000000000000000",55390 => "0000000000000000",
55391 => "0000000000000000",55392 => "0000000000000000",
55393 => "0000000000000000",55394 => "0000000000000000",
55395 => "0000000000000000",55396 => "0000000000000000",
55397 => "0000000000000000",55398 => "0000000000000000",
55399 => "0000000000000000",55400 => "0000000000000000",
55401 => "0000000000000000",55402 => "0000000000000000",
55403 => "0000000000000000",55404 => "0000000000000000",
55405 => "0000000000000000",55406 => "0000000000000000",
55407 => "0000000000000000",55408 => "0000000000000000",
55409 => "0000000000000000",55410 => "0000000000000000",
55411 => "0000000000000000",55412 => "0000000000000000",
55413 => "0000000000000000",55414 => "0000000000000000",
55415 => "0000000000000000",55416 => "0000000000000000",
55417 => "0000000000000000",55418 => "0000000000000000",
55419 => "0000000000000000",55420 => "0000000000000000",
55421 => "0000000000000000",55422 => "0000000000000000",
55423 => "0000000000000000",55424 => "0000000000000000",
55425 => "0000000000000000",55426 => "0000000000000000",
55427 => "0000000000000000",55428 => "0000000000000000",
55429 => "0000000000000000",55430 => "0000000000000000",
55431 => "0000000000000000",55432 => "0000000000000000",
55433 => "0000000000000000",55434 => "0000000000000000",
55435 => "0000000000000000",55436 => "0000000000000000",
55437 => "0000000000000000",55438 => "0000000000000000",
55439 => "0000000000000000",55440 => "0000000000000000",
55441 => "0000000000000000",55442 => "0000000000000000",
55443 => "0000000000000000",55444 => "0000000000000000",
55445 => "0000000000000000",55446 => "0000000000000000",
55447 => "0000000000000000",55448 => "0000000000000000",
55449 => "0000000000000000",55450 => "0000000000000000",
55451 => "0000000000000000",55452 => "0000000000000000",
55453 => "0000000000000000",55454 => "0000000000000000",
55455 => "0000000000000000",55456 => "0000000000000000",
55457 => "0000000000000000",55458 => "0000000000000000",
55459 => "0000000000000000",55460 => "0000000000000000",
55461 => "0000000000000000",55462 => "0000000000000000",
55463 => "0000000000000000",55464 => "0000000000000000",
55465 => "0000000000000000",55466 => "0000000000000000",
55467 => "0000000000000000",55468 => "0000000000000000",
55469 => "0000000000000000",55470 => "0000000000000000",
55471 => "0000000000000000",55472 => "0000000000000000",
55473 => "0000000000000000",55474 => "0000000000000000",
55475 => "0000000000000000",55476 => "0000000000000000",
55477 => "0000000000000000",55478 => "0000000000000000",
55479 => "0000000000000000",55480 => "0000000000000000",
55481 => "0000000000000000",55482 => "0000000000000000",
55483 => "0000000000000000",55484 => "0000000000000000",
55485 => "0000000000000000",55486 => "0000000000000000",
55487 => "0000000000000000",55488 => "0000000000000000",
55489 => "0000000000000000",55490 => "0000000000000000",
55491 => "0000000000000000",55492 => "0000000000000000",
55493 => "0000000000000000",55494 => "0000000000000000",
55495 => "0000000000000000",55496 => "0000000000000000",
55497 => "0000000000000000",55498 => "0000000000000000",
55499 => "0000000000000000",55500 => "0000000000000000",
55501 => "0000000000000000",55502 => "0000000000000000",
55503 => "0000000000000000",55504 => "0000000000000000",
55505 => "0000000000000000",55506 => "0000000000000000",
55507 => "0000000000000000",55508 => "0000000000000000",
55509 => "0000000000000000",55510 => "0000000000000000",
55511 => "0000000000000000",55512 => "0000000000000000",
55513 => "0000000000000000",55514 => "0000000000000000",
55515 => "0000000000000000",55516 => "0000000000000000",
55517 => "0000000000000000",55518 => "0000000000000000",
55519 => "0000000000000000",55520 => "0000000000000000",
55521 => "0000000000000000",55522 => "0000000000000000",
55523 => "0000000000000000",55524 => "0000000000000000",
55525 => "0000000000000000",55526 => "0000000000000000",
55527 => "0000000000000000",55528 => "0000000000000000",
55529 => "0000000000000000",55530 => "0000000000000000",
55531 => "0000000000000000",55532 => "0000000000000000",
55533 => "0000000000000000",55534 => "0000000000000000",
55535 => "0000000000000000",55536 => "0000000000000000",
55537 => "0000000000000000",55538 => "0000000000000000",
55539 => "0000000000000000",55540 => "0000000000000000",
55541 => "0000000000000000",55542 => "0000000000000000",
55543 => "0000000000000000",55544 => "0000000000000000",
55545 => "0000000000000000",55546 => "0000000000000000",
55547 => "0000000000000000",55548 => "0000000000000000",
55549 => "0000000000000000",55550 => "0000000000000000",
55551 => "0000000000000000",55552 => "0000000000000000",
55553 => "0000000000000000",55554 => "0000000000000000",
55555 => "0000000000000000",55556 => "0000000000000000",
55557 => "0000000000000000",55558 => "0000000000000000",
55559 => "0000000000000000",55560 => "0000000000000000",
55561 => "0000000000000000",55562 => "0000000000000000",
55563 => "0000000000000000",55564 => "0000000000000000",
55565 => "0000000000000000",55566 => "0000000000000000",
55567 => "0000000000000000",55568 => "0000000000000000",
55569 => "0000000000000000",55570 => "0000000000000000",
55571 => "0000000000000000",55572 => "0000000000000000",
55573 => "0000000000000000",55574 => "0000000000000000",
55575 => "0000000000000000",55576 => "0000000000000000",
55577 => "0000000000000000",55578 => "0000000000000000",
55579 => "0000000000000000",55580 => "0000000000000000",
55581 => "0000000000000000",55582 => "0000000000000000",
55583 => "0000000000000000",55584 => "0000000000000000",
55585 => "0000000000000000",55586 => "0000000000000000",
55587 => "0000000000000000",55588 => "0000000000000000",
55589 => "0000000000000000",55590 => "0000000000000000",
55591 => "0000000000000000",55592 => "0000000000000000",
55593 => "0000000000000000",55594 => "0000000000000000",
55595 => "0000000000000000",55596 => "0000000000000000",
55597 => "0000000000000000",55598 => "0000000000000000",
55599 => "0000000000000000",55600 => "0000000000000000",
55601 => "0000000000000000",55602 => "0000000000000000",
55603 => "0000000000000000",55604 => "0000000000000000",
55605 => "0000000000000000",55606 => "0000000000000000",
55607 => "0000000000000000",55608 => "0000000000000000",
55609 => "0000000000000000",55610 => "0000000000000000",
55611 => "0000000000000000",55612 => "0000000000000000",
55613 => "0000000000000000",55614 => "0000000000000000",
55615 => "0000000000000000",55616 => "0000000000000000",
55617 => "0000000000000000",55618 => "0000000000000000",
55619 => "0000000000000000",55620 => "0000000000000000",
55621 => "0000000000000000",55622 => "0000000000000000",
55623 => "0000000000000000",55624 => "0000000000000000",
55625 => "0000000000000000",55626 => "0000000000000000",
55627 => "0000000000000000",55628 => "0000000000000000",
55629 => "0000000000000000",55630 => "0000000000000000",
55631 => "0000000000000000",55632 => "0000000000000000",
55633 => "0000000000000000",55634 => "0000000000000000",
55635 => "0000000000000000",55636 => "0000000000000000",
55637 => "0000000000000000",55638 => "0000000000000000",
55639 => "0000000000000000",55640 => "0000000000000000",
55641 => "0000000000000000",55642 => "0000000000000000",
55643 => "0000000000000000",55644 => "0000000000000000",
55645 => "0000000000000000",55646 => "0000000000000000",
55647 => "0000000000000000",55648 => "0000000000000000",
55649 => "0000000000000000",55650 => "0000000000000000",
55651 => "0000000000000000",55652 => "0000000000000000",
55653 => "0000000000000000",55654 => "0000000000000000",
55655 => "0000000000000000",55656 => "0000000000000000",
55657 => "0000000000000000",55658 => "0000000000000000",
55659 => "0000000000000000",55660 => "0000000000000000",
55661 => "0000000000000000",55662 => "0000000000000000",
55663 => "0000000000000000",55664 => "0000000000000000",
55665 => "0000000000000000",55666 => "0000000000000000",
55667 => "0000000000000000",55668 => "0000000000000000",
55669 => "0000000000000000",55670 => "0000000000000000",
55671 => "0000000000000000",55672 => "0000000000000000",
55673 => "0000000000000000",55674 => "0000000000000000",
55675 => "0000000000000000",55676 => "0000000000000000",
55677 => "0000000000000000",55678 => "0000000000000000",
55679 => "0000000000000000",55680 => "0000000000000000",
55681 => "0000000000000000",55682 => "0000000000000000",
55683 => "0000000000000000",55684 => "0000000000000000",
55685 => "0000000000000000",55686 => "0000000000000000",
55687 => "0000000000000000",55688 => "0000000000000000",
55689 => "0000000000000000",55690 => "0000000000000000",
55691 => "0000000000000000",55692 => "0000000000000000",
55693 => "0000000000000000",55694 => "0000000000000000",
55695 => "0000000000000000",55696 => "0000000000000000",
55697 => "0000000000000000",55698 => "0000000000000000",
55699 => "0000000000000000",55700 => "0000000000000000",
55701 => "0000000000000000",55702 => "0000000000000000",
55703 => "0000000000000000",55704 => "0000000000000000",
55705 => "0000000000000000",55706 => "0000000000000000",
55707 => "0000000000000000",55708 => "0000000000000000",
55709 => "0000000000000000",55710 => "0000000000000000",
55711 => "0000000000000000",55712 => "0000000000000000",
55713 => "0000000000000000",55714 => "0000000000000000",
55715 => "0000000000000000",55716 => "0000000000000000",
55717 => "0000000000000000",55718 => "0000000000000000",
55719 => "0000000000000000",55720 => "0000000000000000",
55721 => "0000000000000000",55722 => "0000000000000000",
55723 => "0000000000000000",55724 => "0000000000000000",
55725 => "0000000000000000",55726 => "0000000000000000",
55727 => "0000000000000000",55728 => "0000000000000000",
55729 => "0000000000000000",55730 => "0000000000000000",
55731 => "0000000000000000",55732 => "0000000000000000",
55733 => "0000000000000000",55734 => "0000000000000000",
55735 => "0000000000000000",55736 => "0000000000000000",
55737 => "0000000000000000",55738 => "0000000000000000",
55739 => "0000000000000000",55740 => "0000000000000000",
55741 => "0000000000000000",55742 => "0000000000000000",
55743 => "0000000000000000",55744 => "0000000000000000",
55745 => "0000000000000000",55746 => "0000000000000000",
55747 => "0000000000000000",55748 => "0000000000000000",
55749 => "0000000000000000",55750 => "0000000000000000",
55751 => "0000000000000000",55752 => "0000000000000000",
55753 => "0000000000000000",55754 => "0000000000000000",
55755 => "0000000000000000",55756 => "0000000000000000",
55757 => "0000000000000000",55758 => "0000000000000000",
55759 => "0000000000000000",55760 => "0000000000000000",
55761 => "0000000000000000",55762 => "0000000000000000",
55763 => "0000000000000000",55764 => "0000000000000000",
55765 => "0000000000000000",55766 => "0000000000000000",
55767 => "0000000000000000",55768 => "0000000000000000",
55769 => "0000000000000000",55770 => "0000000000000000",
55771 => "0000000000000000",55772 => "0000000000000000",
55773 => "0000000000000000",55774 => "0000000000000000",
55775 => "0000000000000000",55776 => "0000000000000000",
55777 => "0000000000000000",55778 => "0000000000000000",
55779 => "0000000000000000",55780 => "0000000000000000",
55781 => "0000000000000000",55782 => "0000000000000000",
55783 => "0000000000000000",55784 => "0000000000000000",
55785 => "0000000000000000",55786 => "0000000000000000",
55787 => "0000000000000000",55788 => "0000000000000000",
55789 => "0000000000000000",55790 => "0000000000000000",
55791 => "0000000000000000",55792 => "0000000000000000",
55793 => "0000000000000000",55794 => "0000000000000000",
55795 => "0000000000000000",55796 => "0000000000000000",
55797 => "0000000000000000",55798 => "0000000000000000",
55799 => "0000000000000000",55800 => "0000000000000000",
55801 => "0000000000000000",55802 => "0000000000000000",
55803 => "0000000000000000",55804 => "0000000000000000",
55805 => "0000000000000000",55806 => "0000000000000000",
55807 => "0000000000000000",55808 => "0000000000000000",
55809 => "0000000000000000",55810 => "0000000000000000",
55811 => "0000000000000000",55812 => "0000000000000000",
55813 => "0000000000000000",55814 => "0000000000000000",
55815 => "0000000000000000",55816 => "0000000000000000",
55817 => "0000000000000000",55818 => "0000000000000000",
55819 => "0000000000000000",55820 => "0000000000000000",
55821 => "0000000000000000",55822 => "0000000000000000",
55823 => "0000000000000000",55824 => "0000000000000000",
55825 => "0000000000000000",55826 => "0000000000000000",
55827 => "0000000000000000",55828 => "0000000000000000",
55829 => "0000000000000000",55830 => "0000000000000000",
55831 => "0000000000000000",55832 => "0000000000000000",
55833 => "0000000000000000",55834 => "0000000000000000",
55835 => "0000000000000000",55836 => "0000000000000000",
55837 => "0000000000000000",55838 => "0000000000000000",
55839 => "0000000000000000",55840 => "0000000000000000",
55841 => "0000000000000000",55842 => "0000000000000000",
55843 => "0000000000000000",55844 => "0000000000000000",
55845 => "0000000000000000",55846 => "0000000000000000",
55847 => "0000000000000000",55848 => "0000000000000000",
55849 => "0000000000000000",55850 => "0000000000000000",
55851 => "0000000000000000",55852 => "0000000000000000",
55853 => "0000000000000000",55854 => "0000000000000000",
55855 => "0000000000000000",55856 => "0000000000000000",
55857 => "0000000000000000",55858 => "0000000000000000",
55859 => "0000000000000000",55860 => "0000000000000000",
55861 => "0000000000000000",55862 => "0000000000000000",
55863 => "0000000000000000",55864 => "0000000000000000",
55865 => "0000000000000000",55866 => "0000000000000000",
55867 => "0000000000000000",55868 => "0000000000000000",
55869 => "0000000000000000",55870 => "0000000000000000",
55871 => "0000000000000000",55872 => "0000000000000000",
55873 => "0000000000000000",55874 => "0000000000000000",
55875 => "0000000000000000",55876 => "0000000000000000",
55877 => "0000000000000000",55878 => "0000000000000000",
55879 => "0000000000000000",55880 => "0000000000000000",
55881 => "0000000000000000",55882 => "0000000000000000",
55883 => "0000000000000000",55884 => "0000000000000000",
55885 => "0000000000000000",55886 => "0000000000000000",
55887 => "0000000000000000",55888 => "0000000000000000",
55889 => "0000000000000000",55890 => "0000000000000000",
55891 => "0000000000000000",55892 => "0000000000000000",
55893 => "0000000000000000",55894 => "0000000000000000",
55895 => "0000000000000000",55896 => "0000000000000000",
55897 => "0000000000000000",55898 => "0000000000000000",
55899 => "0000000000000000",55900 => "0000000000000000",
55901 => "0000000000000000",55902 => "0000000000000000",
55903 => "0000000000000000",55904 => "0000000000000000",
55905 => "0000000000000000",55906 => "0000000000000000",
55907 => "0000000000000000",55908 => "0000000000000000",
55909 => "0000000000000000",55910 => "0000000000000000",
55911 => "0000000000000000",55912 => "0000000000000000",
55913 => "0000000000000000",55914 => "0000000000000000",
55915 => "0000000000000000",55916 => "0000000000000000",
55917 => "0000000000000000",55918 => "0000000000000000",
55919 => "0000000000000000",55920 => "0000000000000000",
55921 => "0000000000000000",55922 => "0000000000000000",
55923 => "0000000000000000",55924 => "0000000000000000",
55925 => "0000000000000000",55926 => "0000000000000000",
55927 => "0000000000000000",55928 => "0000000000000000",
55929 => "0000000000000000",55930 => "0000000000000000",
55931 => "0000000000000000",55932 => "0000000000000000",
55933 => "0000000000000000",55934 => "0000000000000000",
55935 => "0000000000000000",55936 => "0000000000000000",
55937 => "0000000000000000",55938 => "0000000000000000",
55939 => "0000000000000000",55940 => "0000000000000000",
55941 => "0000000000000000",55942 => "0000000000000000",
55943 => "0000000000000000",55944 => "0000000000000000",
55945 => "0000000000000000",55946 => "0000000000000000",
55947 => "0000000000000000",55948 => "0000000000000000",
55949 => "0000000000000000",55950 => "0000000000000000",
55951 => "0000000000000000",55952 => "0000000000000000",
55953 => "0000000000000000",55954 => "0000000000000000",
55955 => "0000000000000000",55956 => "0000000000000000",
55957 => "0000000000000000",55958 => "0000000000000000",
55959 => "0000000000000000",55960 => "0000000000000000",
55961 => "0000000000000000",55962 => "0000000000000000",
55963 => "0000000000000000",55964 => "0000000000000000",
55965 => "0000000000000000",55966 => "0000000000000000",
55967 => "0000000000000000",55968 => "0000000000000000",
55969 => "0000000000000000",55970 => "0000000000000000",
55971 => "0000000000000000",55972 => "0000000000000000",
55973 => "0000000000000000",55974 => "0000000000000000",
55975 => "0000000000000000",55976 => "0000000000000000",
55977 => "0000000000000000",55978 => "0000000000000000",
55979 => "0000000000000000",55980 => "0000000000000000",
55981 => "0000000000000000",55982 => "0000000000000000",
55983 => "0000000000000000",55984 => "0000000000000000",
55985 => "0000000000000000",55986 => "0000000000000000",
55987 => "0000000000000000",55988 => "0000000000000000",
55989 => "0000000000000000",55990 => "0000000000000000",
55991 => "0000000000000000",55992 => "0000000000000000",
55993 => "0000000000000000",55994 => "0000000000000000",
55995 => "0000000000000000",55996 => "0000000000000000",
55997 => "0000000000000000",55998 => "0000000000000000",
55999 => "0000000000000000",56000 => "0000000000000000",
56001 => "0000000000000000",56002 => "0000000000000000",
56003 => "0000000000000000",56004 => "0000000000000000",
56005 => "0000000000000000",56006 => "0000000000000000",
56007 => "0000000000000000",56008 => "0000000000000000",
56009 => "0000000000000000",56010 => "0000000000000000",
56011 => "0000000000000000",56012 => "0000000000000000",
56013 => "0000000000000000",56014 => "0000000000000000",
56015 => "0000000000000000",56016 => "0000000000000000",
56017 => "0000000000000000",56018 => "0000000000000000",
56019 => "0000000000000000",56020 => "0000000000000000",
56021 => "0000000000000000",56022 => "0000000000000000",
56023 => "0000000000000000",56024 => "0000000000000000",
56025 => "0000000000000000",56026 => "0000000000000000",
56027 => "0000000000000000",56028 => "0000000000000000",
56029 => "0000000000000000",56030 => "0000000000000000",
56031 => "0000000000000000",56032 => "0000000000000000",
56033 => "0000000000000000",56034 => "0000000000000000",
56035 => "0000000000000000",56036 => "0000000000000000",
56037 => "0000000000000000",56038 => "0000000000000000",
56039 => "0000000000000000",56040 => "0000000000000000",
56041 => "0000000000000000",56042 => "0000000000000000",
56043 => "0000000000000000",56044 => "0000000000000000",
56045 => "0000000000000000",56046 => "0000000000000000",
56047 => "0000000000000000",56048 => "0000000000000000",
56049 => "0000000000000000",56050 => "0000000000000000",
56051 => "0000000000000000",56052 => "0000000000000000",
56053 => "0000000000000000",56054 => "0000000000000000",
56055 => "0000000000000000",56056 => "0000000000000000",
56057 => "0000000000000000",56058 => "0000000000000000",
56059 => "0000000000000000",56060 => "0000000000000000",
56061 => "0000000000000000",56062 => "0000000000000000",
56063 => "0000000000000000",56064 => "0000000000000000",
56065 => "0000000000000000",56066 => "0000000000000000",
56067 => "0000000000000000",56068 => "0000000000000000",
56069 => "0000000000000000",56070 => "0000000000000000",
56071 => "0000000000000000",56072 => "0000000000000000",
56073 => "0000000000000000",56074 => "0000000000000000",
56075 => "0000000000000000",56076 => "0000000000000000",
56077 => "0000000000000000",56078 => "0000000000000000",
56079 => "0000000000000000",56080 => "0000000000000000",
56081 => "0000000000000000",56082 => "0000000000000000",
56083 => "0000000000000000",56084 => "0000000000000000",
56085 => "0000000000000000",56086 => "0000000000000000",
56087 => "0000000000000000",56088 => "0000000000000000",
56089 => "0000000000000000",56090 => "0000000000000000",
56091 => "0000000000000000",56092 => "0000000000000000",
56093 => "0000000000000000",56094 => "0000000000000000",
56095 => "0000000000000000",56096 => "0000000000000000",
56097 => "0000000000000000",56098 => "0000000000000000",
56099 => "0000000000000000",56100 => "0000000000000000",
56101 => "0000000000000000",56102 => "0000000000000000",
56103 => "0000000000000000",56104 => "0000000000000000",
56105 => "0000000000000000",56106 => "0000000000000000",
56107 => "0000000000000000",56108 => "0000000000000000",
56109 => "0000000000000000",56110 => "0000000000000000",
56111 => "0000000000000000",56112 => "0000000000000000",
56113 => "0000000000000000",56114 => "0000000000000000",
56115 => "0000000000000000",56116 => "0000000000000000",
56117 => "0000000000000000",56118 => "0000000000000000",
56119 => "0000000000000000",56120 => "0000000000000000",
56121 => "0000000000000000",56122 => "0000000000000000",
56123 => "0000000000000000",56124 => "0000000000000000",
56125 => "0000000000000000",56126 => "0000000000000000",
56127 => "0000000000000000",56128 => "0000000000000000",
56129 => "0000000000000000",56130 => "0000000000000000",
56131 => "0000000000000000",56132 => "0000000000000000",
56133 => "0000000000000000",56134 => "0000000000000000",
56135 => "0000000000000000",56136 => "0000000000000000",
56137 => "0000000000000000",56138 => "0000000000000000",
56139 => "0000000000000000",56140 => "0000000000000000",
56141 => "0000000000000000",56142 => "0000000000000000",
56143 => "0000000000000000",56144 => "0000000000000000",
56145 => "0000000000000000",56146 => "0000000000000000",
56147 => "0000000000000000",56148 => "0000000000000000",
56149 => "0000000000000000",56150 => "0000000000000000",
56151 => "0000000000000000",56152 => "0000000000000000",
56153 => "0000000000000000",56154 => "0000000000000000",
56155 => "0000000000000000",56156 => "0000000000000000",
56157 => "0000000000000000",56158 => "0000000000000000",
56159 => "0000000000000000",56160 => "0000000000000000",
56161 => "0000000000000000",56162 => "0000000000000000",
56163 => "0000000000000000",56164 => "0000000000000000",
56165 => "0000000000000000",56166 => "0000000000000000",
56167 => "0000000000000000",56168 => "0000000000000000",
56169 => "0000000000000000",56170 => "0000000000000000",
56171 => "0000000000000000",56172 => "0000000000000000",
56173 => "0000000000000000",56174 => "0000000000000000",
56175 => "0000000000000000",56176 => "0000000000000000",
56177 => "0000000000000000",56178 => "0000000000000000",
56179 => "0000000000000000",56180 => "0000000000000000",
56181 => "0000000000000000",56182 => "0000000000000000",
56183 => "0000000000000000",56184 => "0000000000000000",
56185 => "0000000000000000",56186 => "0000000000000000",
56187 => "0000000000000000",56188 => "0000000000000000",
56189 => "0000000000000000",56190 => "0000000000000000",
56191 => "0000000000000000",56192 => "0000000000000000",
56193 => "0000000000000000",56194 => "0000000000000000",
56195 => "0000000000000000",56196 => "0000000000000000",
56197 => "0000000000000000",56198 => "0000000000000000",
56199 => "0000000000000000",56200 => "0000000000000000",
56201 => "0000000000000000",56202 => "0000000000000000",
56203 => "0000000000000000",56204 => "0000000000000000",
56205 => "0000000000000000",56206 => "0000000000000000",
56207 => "0000000000000000",56208 => "0000000000000000",
56209 => "0000000000000000",56210 => "0000000000000000",
56211 => "0000000000000000",56212 => "0000000000000000",
56213 => "0000000000000000",56214 => "0000000000000000",
56215 => "0000000000000000",56216 => "0000000000000000",
56217 => "0000000000000000",56218 => "0000000000000000",
56219 => "0000000000000000",56220 => "0000000000000000",
56221 => "0000000000000000",56222 => "0000000000000000",
56223 => "0000000000000000",56224 => "0000000000000000",
56225 => "0000000000000000",56226 => "0000000000000000",
56227 => "0000000000000000",56228 => "0000000000000000",
56229 => "0000000000000000",56230 => "0000000000000000",
56231 => "0000000000000000",56232 => "0000000000000000",
56233 => "0000000000000000",56234 => "0000000000000000",
56235 => "0000000000000000",56236 => "0000000000000000",
56237 => "0000000000000000",56238 => "0000000000000000",
56239 => "0000000000000000",56240 => "0000000000000000",
56241 => "0000000000000000",56242 => "0000000000000000",
56243 => "0000000000000000",56244 => "0000000000000000",
56245 => "0000000000000000",56246 => "0000000000000000",
56247 => "0000000000000000",56248 => "0000000000000000",
56249 => "0000000000000000",56250 => "0000000000000000",
56251 => "0000000000000000",56252 => "0000000000000000",
56253 => "0000000000000000",56254 => "0000000000000000",
56255 => "0000000000000000",56256 => "0000000000000000",
56257 => "0000000000000000",56258 => "0000000000000000",
56259 => "0000000000000000",56260 => "0000000000000000",
56261 => "0000000000000000",56262 => "0000000000000000",
56263 => "0000000000000000",56264 => "0000000000000000",
56265 => "0000000000000000",56266 => "0000000000000000",
56267 => "0000000000000000",56268 => "0000000000000000",
56269 => "0000000000000000",56270 => "0000000000000000",
56271 => "0000000000000000",56272 => "0000000000000000",
56273 => "0000000000000000",56274 => "0000000000000000",
56275 => "0000000000000000",56276 => "0000000000000000",
56277 => "0000000000000000",56278 => "0000000000000000",
56279 => "0000000000000000",56280 => "0000000000000000",
56281 => "0000000000000000",56282 => "0000000000000000",
56283 => "0000000000000000",56284 => "0000000000000000",
56285 => "0000000000000000",56286 => "0000000000000000",
56287 => "0000000000000000",56288 => "0000000000000000",
56289 => "0000000000000000",56290 => "0000000000000000",
56291 => "0000000000000000",56292 => "0000000000000000",
56293 => "0000000000000000",56294 => "0000000000000000",
56295 => "0000000000000000",56296 => "0000000000000000",
56297 => "0000000000000000",56298 => "0000000000000000",
56299 => "0000000000000000",56300 => "0000000000000000",
56301 => "0000000000000000",56302 => "0000000000000000",
56303 => "0000000000000000",56304 => "0000000000000000",
56305 => "0000000000000000",56306 => "0000000000000000",
56307 => "0000000000000000",56308 => "0000000000000000",
56309 => "0000000000000000",56310 => "0000000000000000",
56311 => "0000000000000000",56312 => "0000000000000000",
56313 => "0000000000000000",56314 => "0000000000000000",
56315 => "0000000000000000",56316 => "0000000000000000",
56317 => "0000000000000000",56318 => "0000000000000000",
56319 => "0000000000000000",56320 => "0000000000000000",
56321 => "0000000000000000",56322 => "0000000000000000",
56323 => "0000000000000000",56324 => "0000000000000000",
56325 => "0000000000000000",56326 => "0000000000000000",
56327 => "0000000000000000",56328 => "0000000000000000",
56329 => "0000000000000000",56330 => "0000000000000000",
56331 => "0000000000000000",56332 => "0000000000000000",
56333 => "0000000000000000",56334 => "0000000000000000",
56335 => "0000000000000000",56336 => "0000000000000000",
56337 => "0000000000000000",56338 => "0000000000000000",
56339 => "0000000000000000",56340 => "0000000000000000",
56341 => "0000000000000000",56342 => "0000000000000000",
56343 => "0000000000000000",56344 => "0000000000000000",
56345 => "0000000000000000",56346 => "0000000000000000",
56347 => "0000000000000000",56348 => "0000000000000000",
56349 => "0000000000000000",56350 => "0000000000000000",
56351 => "0000000000000000",56352 => "0000000000000000",
56353 => "0000000000000000",56354 => "0000000000000000",
56355 => "0000000000000000",56356 => "0000000000000000",
56357 => "0000000000000000",56358 => "0000000000000000",
56359 => "0000000000000000",56360 => "0000000000000000",
56361 => "0000000000000000",56362 => "0000000000000000",
56363 => "0000000000000000",56364 => "0000000000000000",
56365 => "0000000000000000",56366 => "0000000000000000",
56367 => "0000000000000000",56368 => "0000000000000000",
56369 => "0000000000000000",56370 => "0000000000000000",
56371 => "0000000000000000",56372 => "0000000000000000",
56373 => "0000000000000000",56374 => "0000000000000000",
56375 => "0000000000000000",56376 => "0000000000000000",
56377 => "0000000000000000",56378 => "0000000000000000",
56379 => "0000000000000000",56380 => "0000000000000000",
56381 => "0000000000000000",56382 => "0000000000000000",
56383 => "0000000000000000",56384 => "0000000000000000",
56385 => "0000000000000000",56386 => "0000000000000000",
56387 => "0000000000000000",56388 => "0000000000000000",
56389 => "0000000000000000",56390 => "0000000000000000",
56391 => "0000000000000000",56392 => "0000000000000000",
56393 => "0000000000000000",56394 => "0000000000000000",
56395 => "0000000000000000",56396 => "0000000000000000",
56397 => "0000000000000000",56398 => "0000000000000000",
56399 => "0000000000000000",56400 => "0000000000000000",
56401 => "0000000000000000",56402 => "0000000000000000",
56403 => "0000000000000000",56404 => "0000000000000000",
56405 => "0000000000000000",56406 => "0000000000000000",
56407 => "0000000000000000",56408 => "0000000000000000",
56409 => "0000000000000000",56410 => "0000000000000000",
56411 => "0000000000000000",56412 => "0000000000000000",
56413 => "0000000000000000",56414 => "0000000000000000",
56415 => "0000000000000000",56416 => "0000000000000000",
56417 => "0000000000000000",56418 => "0000000000000000",
56419 => "0000000000000000",56420 => "0000000000000000",
56421 => "0000000000000000",56422 => "0000000000000000",
56423 => "0000000000000000",56424 => "0000000000000000",
56425 => "0000000000000000",56426 => "0000000000000000",
56427 => "0000000000000000",56428 => "0000000000000000",
56429 => "0000000000000000",56430 => "0000000000000000",
56431 => "0000000000000000",56432 => "0000000000000000",
56433 => "0000000000000000",56434 => "0000000000000000",
56435 => "0000000000000000",56436 => "0000000000000000",
56437 => "0000000000000000",56438 => "0000000000000000",
56439 => "0000000000000000",56440 => "0000000000000000",
56441 => "0000000000000000",56442 => "0000000000000000",
56443 => "0000000000000000",56444 => "0000000000000000",
56445 => "0000000000000000",56446 => "0000000000000000",
56447 => "0000000000000000",56448 => "0000000000000000",
56449 => "0000000000000000",56450 => "0000000000000000",
56451 => "0000000000000000",56452 => "0000000000000000",
56453 => "0000000000000000",56454 => "0000000000000000",
56455 => "0000000000000000",56456 => "0000000000000000",
56457 => "0000000000000000",56458 => "0000000000000000",
56459 => "0000000000000000",56460 => "0000000000000000",
56461 => "0000000000000000",56462 => "0000000000000000",
56463 => "0000000000000000",56464 => "0000000000000000",
56465 => "0000000000000000",56466 => "0000000000000000",
56467 => "0000000000000000",56468 => "0000000000000000",
56469 => "0000000000000000",56470 => "0000000000000000",
56471 => "0000000000000000",56472 => "0000000000000000",
56473 => "0000000000000000",56474 => "0000000000000000",
56475 => "0000000000000000",56476 => "0000000000000000",
56477 => "0000000000000000",56478 => "0000000000000000",
56479 => "0000000000000000",56480 => "0000000000000000",
56481 => "0000000000000000",56482 => "0000000000000000",
56483 => "0000000000000000",56484 => "0000000000000000",
56485 => "0000000000000000",56486 => "0000000000000000",
56487 => "0000000000000000",56488 => "0000000000000000",
56489 => "0000000000000000",56490 => "0000000000000000",
56491 => "0000000000000000",56492 => "0000000000000000",
56493 => "0000000000000000",56494 => "0000000000000000",
56495 => "0000000000000000",56496 => "0000000000000000",
56497 => "0000000000000000",56498 => "0000000000000000",
56499 => "0000000000000000",56500 => "0000000000000000",
56501 => "0000000000000000",56502 => "0000000000000000",
56503 => "0000000000000000",56504 => "0000000000000000",
56505 => "0000000000000000",56506 => "0000000000000000",
56507 => "0000000000000000",56508 => "0000000000000000",
56509 => "0000000000000000",56510 => "0000000000000000",
56511 => "0000000000000000",56512 => "0000000000000000",
56513 => "0000000000000000",56514 => "0000000000000000",
56515 => "0000000000000000",56516 => "0000000000000000",
56517 => "0000000000000000",56518 => "0000000000000000",
56519 => "0000000000000000",56520 => "0000000000000000",
56521 => "0000000000000000",56522 => "0000000000000000",
56523 => "0000000000000000",56524 => "0000000000000000",
56525 => "0000000000000000",56526 => "0000000000000000",
56527 => "0000000000000000",56528 => "0000000000000000",
56529 => "0000000000000000",56530 => "0000000000000000",
56531 => "0000000000000000",56532 => "0000000000000000",
56533 => "0000000000000000",56534 => "0000000000000000",
56535 => "0000000000000000",56536 => "0000000000000000",
56537 => "0000000000000000",56538 => "0000000000000000",
56539 => "0000000000000000",56540 => "0000000000000000",
56541 => "0000000000000000",56542 => "0000000000000000",
56543 => "0000000000000000",56544 => "0000000000000000",
56545 => "0000000000000000",56546 => "0000000000000000",
56547 => "0000000000000000",56548 => "0000000000000000",
56549 => "0000000000000000",56550 => "0000000000000000",
56551 => "0000000000000000",56552 => "0000000000000000",
56553 => "0000000000000000",56554 => "0000000000000000",
56555 => "0000000000000000",56556 => "0000000000000000",
56557 => "0000000000000000",56558 => "0000000000000000",
56559 => "0000000000000000",56560 => "0000000000000000",
56561 => "0000000000000000",56562 => "0000000000000000",
56563 => "0000000000000000",56564 => "0000000000000000",
56565 => "0000000000000000",56566 => "0000000000000000",
56567 => "0000000000000000",56568 => "0000000000000000",
56569 => "0000000000000000",56570 => "0000000000000000",
56571 => "0000000000000000",56572 => "0000000000000000",
56573 => "0000000000000000",56574 => "0000000000000000",
56575 => "0000000000000000",56576 => "0000000000000000",
56577 => "0000000000000000",56578 => "0000000000000000",
56579 => "0000000000000000",56580 => "0000000000000000",
56581 => "0000000000000000",56582 => "0000000000000000",
56583 => "0000000000000000",56584 => "0000000000000000",
56585 => "0000000000000000",56586 => "0000000000000000",
56587 => "0000000000000000",56588 => "0000000000000000",
56589 => "0000000000000000",56590 => "0000000000000000",
56591 => "0000000000000000",56592 => "0000000000000000",
56593 => "0000000000000000",56594 => "0000000000000000",
56595 => "0000000000000000",56596 => "0000000000000000",
56597 => "0000000000000000",56598 => "0000000000000000",
56599 => "0000000000000000",56600 => "0000000000000000",
56601 => "0000000000000000",56602 => "0000000000000000",
56603 => "0000000000000000",56604 => "0000000000000000",
56605 => "0000000000000000",56606 => "0000000000000000",
56607 => "0000000000000000",56608 => "0000000000000000",
56609 => "0000000000000000",56610 => "0000000000000000",
56611 => "0000000000000000",56612 => "0000000000000000",
56613 => "0000000000000000",56614 => "0000000000000000",
56615 => "0000000000000000",56616 => "0000000000000000",
56617 => "0000000000000000",56618 => "0000000000000000",
56619 => "0000000000000000",56620 => "0000000000000000",
56621 => "0000000000000000",56622 => "0000000000000000",
56623 => "0000000000000000",56624 => "0000000000000000",
56625 => "0000000000000000",56626 => "0000000000000000",
56627 => "0000000000000000",56628 => "0000000000000000",
56629 => "0000000000000000",56630 => "0000000000000000",
56631 => "0000000000000000",56632 => "0000000000000000",
56633 => "0000000000000000",56634 => "0000000000000000",
56635 => "0000000000000000",56636 => "0000000000000000",
56637 => "0000000000000000",56638 => "0000000000000000",
56639 => "0000000000000000",56640 => "0000000000000000",
56641 => "0000000000000000",56642 => "0000000000000000",
56643 => "0000000000000000",56644 => "0000000000000000",
56645 => "0000000000000000",56646 => "0000000000000000",
56647 => "0000000000000000",56648 => "0000000000000000",
56649 => "0000000000000000",56650 => "0000000000000000",
56651 => "0000000000000000",56652 => "0000000000000000",
56653 => "0000000000000000",56654 => "0000000000000000",
56655 => "0000000000000000",56656 => "0000000000000000",
56657 => "0000000000000000",56658 => "0000000000000000",
56659 => "0000000000000000",56660 => "0000000000000000",
56661 => "0000000000000000",56662 => "0000000000000000",
56663 => "0000000000000000",56664 => "0000000000000000",
56665 => "0000000000000000",56666 => "0000000000000000",
56667 => "0000000000000000",56668 => "0000000000000000",
56669 => "0000000000000000",56670 => "0000000000000000",
56671 => "0000000000000000",56672 => "0000000000000000",
56673 => "0000000000000000",56674 => "0000000000000000",
56675 => "0000000000000000",56676 => "0000000000000000",
56677 => "0000000000000000",56678 => "0000000000000000",
56679 => "0000000000000000",56680 => "0000000000000000",
56681 => "0000000000000000",56682 => "0000000000000000",
56683 => "0000000000000000",56684 => "0000000000000000",
56685 => "0000000000000000",56686 => "0000000000000000",
56687 => "0000000000000000",56688 => "0000000000000000",
56689 => "0000000000000000",56690 => "0000000000000000",
56691 => "0000000000000000",56692 => "0000000000000000",
56693 => "0000000000000000",56694 => "0000000000000000",
56695 => "0000000000000000",56696 => "0000000000000000",
56697 => "0000000000000000",56698 => "0000000000000000",
56699 => "0000000000000000",56700 => "0000000000000000",
56701 => "0000000000000000",56702 => "0000000000000000",
56703 => "0000000000000000",56704 => "0000000000000000",
56705 => "0000000000000000",56706 => "0000000000000000",
56707 => "0000000000000000",56708 => "0000000000000000",
56709 => "0000000000000000",56710 => "0000000000000000",
56711 => "0000000000000000",56712 => "0000000000000000",
56713 => "0000000000000000",56714 => "0000000000000000",
56715 => "0000000000000000",56716 => "0000000000000000",
56717 => "0000000000000000",56718 => "0000000000000000",
56719 => "0000000000000000",56720 => "0000000000000000",
56721 => "0000000000000000",56722 => "0000000000000000",
56723 => "0000000000000000",56724 => "0000000000000000",
56725 => "0000000000000000",56726 => "0000000000000000",
56727 => "0000000000000000",56728 => "0000000000000000",
56729 => "0000000000000000",56730 => "0000000000000000",
56731 => "0000000000000000",56732 => "0000000000000000",
56733 => "0000000000000000",56734 => "0000000000000000",
56735 => "0000000000000000",56736 => "0000000000000000",
56737 => "0000000000000000",56738 => "0000000000000000",
56739 => "0000000000000000",56740 => "0000000000000000",
56741 => "0000000000000000",56742 => "0000000000000000",
56743 => "0000000000000000",56744 => "0000000000000000",
56745 => "0000000000000000",56746 => "0000000000000000",
56747 => "0000000000000000",56748 => "0000000000000000",
56749 => "0000000000000000",56750 => "0000000000000000",
56751 => "0000000000000000",56752 => "0000000000000000",
56753 => "0000000000000000",56754 => "0000000000000000",
56755 => "0000000000000000",56756 => "0000000000000000",
56757 => "0000000000000000",56758 => "0000000000000000",
56759 => "0000000000000000",56760 => "0000000000000000",
56761 => "0000000000000000",56762 => "0000000000000000",
56763 => "0000000000000000",56764 => "0000000000000000",
56765 => "0000000000000000",56766 => "0000000000000000",
56767 => "0000000000000000",56768 => "0000000000000000",
56769 => "0000000000000000",56770 => "0000000000000000",
56771 => "0000000000000000",56772 => "0000000000000000",
56773 => "0000000000000000",56774 => "0000000000000000",
56775 => "0000000000000000",56776 => "0000000000000000",
56777 => "0000000000000000",56778 => "0000000000000000",
56779 => "0000000000000000",56780 => "0000000000000000",
56781 => "0000000000000000",56782 => "0000000000000000",
56783 => "0000000000000000",56784 => "0000000000000000",
56785 => "0000000000000000",56786 => "0000000000000000",
56787 => "0000000000000000",56788 => "0000000000000000",
56789 => "0000000000000000",56790 => "0000000000000000",
56791 => "0000000000000000",56792 => "0000000000000000",
56793 => "0000000000000000",56794 => "0000000000000000",
56795 => "0000000000000000",56796 => "0000000000000000",
56797 => "0000000000000000",56798 => "0000000000000000",
56799 => "0000000000000000",56800 => "0000000000000000",
56801 => "0000000000000000",56802 => "0000000000000000",
56803 => "0000000000000000",56804 => "0000000000000000",
56805 => "0000000000000000",56806 => "0000000000000000",
56807 => "0000000000000000",56808 => "0000000000000000",
56809 => "0000000000000000",56810 => "0000000000000000",
56811 => "0000000000000000",56812 => "0000000000000000",
56813 => "0000000000000000",56814 => "0000000000000000",
56815 => "0000000000000000",56816 => "0000000000000000",
56817 => "0000000000000000",56818 => "0000000000000000",
56819 => "0000000000000000",56820 => "0000000000000000",
56821 => "0000000000000000",56822 => "0000000000000000",
56823 => "0000000000000000",56824 => "0000000000000000",
56825 => "0000000000000000",56826 => "0000000000000000",
56827 => "0000000000000000",56828 => "0000000000000000",
56829 => "0000000000000000",56830 => "0000000000000000",
56831 => "0000000000000000",56832 => "0000000000000000",
56833 => "0000000000000000",56834 => "0000000000000000",
56835 => "0000000000000000",56836 => "0000000000000000",
56837 => "0000000000000000",56838 => "0000000000000000",
56839 => "0000000000000000",56840 => "0000000000000000",
56841 => "0000000000000000",56842 => "0000000000000000",
56843 => "0000000000000000",56844 => "0000000000000000",
56845 => "0000000000000000",56846 => "0000000000000000",
56847 => "0000000000000000",56848 => "0000000000000000",
56849 => "0000000000000000",56850 => "0000000000000000",
56851 => "0000000000000000",56852 => "0000000000000000",
56853 => "0000000000000000",56854 => "0000000000000000",
56855 => "0000000000000000",56856 => "0000000000000000",
56857 => "0000000000000000",56858 => "0000000000000000",
56859 => "0000000000000000",56860 => "0000000000000000",
56861 => "0000000000000000",56862 => "0000000000000000",
56863 => "0000000000000000",56864 => "0000000000000000",
56865 => "0000000000000000",56866 => "0000000000000000",
56867 => "0000000000000000",56868 => "0000000000000000",
56869 => "0000000000000000",56870 => "0000000000000000",
56871 => "0000000000000000",56872 => "0000000000000000",
56873 => "0000000000000000",56874 => "0000000000000000",
56875 => "0000000000000000",56876 => "0000000000000000",
56877 => "0000000000000000",56878 => "0000000000000000",
56879 => "0000000000000000",56880 => "0000000000000000",
56881 => "0000000000000000",56882 => "0000000000000000",
56883 => "0000000000000000",56884 => "0000000000000000",
56885 => "0000000000000000",56886 => "0000000000000000",
56887 => "0000000000000000",56888 => "0000000000000000",
56889 => "0000000000000000",56890 => "0000000000000000",
56891 => "0000000000000000",56892 => "0000000000000000",
56893 => "0000000000000000",56894 => "0000000000000000",
56895 => "0000000000000000",56896 => "0000000000000000",
56897 => "0000000000000000",56898 => "0000000000000000",
56899 => "0000000000000000",56900 => "0000000000000000",
56901 => "0000000000000000",56902 => "0000000000000000",
56903 => "0000000000000000",56904 => "0000000000000000",
56905 => "0000000000000000",56906 => "0000000000000000",
56907 => "0000000000000000",56908 => "0000000000000000",
56909 => "0000000000000000",56910 => "0000000000000000",
56911 => "0000000000000000",56912 => "0000000000000000",
56913 => "0000000000000000",56914 => "0000000000000000",
56915 => "0000000000000000",56916 => "0000000000000000",
56917 => "0000000000000000",56918 => "0000000000000000",
56919 => "0000000000000000",56920 => "0000000000000000",
56921 => "0000000000000000",56922 => "0000000000000000",
56923 => "0000000000000000",56924 => "0000000000000000",
56925 => "0000000000000000",56926 => "0000000000000000",
56927 => "0000000000000000",56928 => "0000000000000000",
56929 => "0000000000000000",56930 => "0000000000000000",
56931 => "0000000000000000",56932 => "0000000000000000",
56933 => "0000000000000000",56934 => "0000000000000000",
56935 => "0000000000000000",56936 => "0000000000000000",
56937 => "0000000000000000",56938 => "0000000000000000",
56939 => "0000000000000000",56940 => "0000000000000000",
56941 => "0000000000000000",56942 => "0000000000000000",
56943 => "0000000000000000",56944 => "0000000000000000",
56945 => "0000000000000000",56946 => "0000000000000000",
56947 => "0000000000000000",56948 => "0000000000000000",
56949 => "0000000000000000",56950 => "0000000000000000",
56951 => "0000000000000000",56952 => "0000000000000000",
56953 => "0000000000000000",56954 => "0000000000000000",
56955 => "0000000000000000",56956 => "0000000000000000",
56957 => "0000000000000000",56958 => "0000000000000000",
56959 => "0000000000000000",56960 => "0000000000000000",
56961 => "0000000000000000",56962 => "0000000000000000",
56963 => "0000000000000000",56964 => "0000000000000000",
56965 => "0000000000000000",56966 => "0000000000000000",
56967 => "0000000000000000",56968 => "0000000000000000",
56969 => "0000000000000000",56970 => "0000000000000000",
56971 => "0000000000000000",56972 => "0000000000000000",
56973 => "0000000000000000",56974 => "0000000000000000",
56975 => "0000000000000000",56976 => "0000000000000000",
56977 => "0000000000000000",56978 => "0000000000000000",
56979 => "0000000000000000",56980 => "0000000000000000",
56981 => "0000000000000000",56982 => "0000000000000000",
56983 => "0000000000000000",56984 => "0000000000000000",
56985 => "0000000000000000",56986 => "0000000000000000",
56987 => "0000000000000000",56988 => "0000000000000000",
56989 => "0000000000000000",56990 => "0000000000000000",
56991 => "0000000000000000",56992 => "0000000000000000",
56993 => "0000000000000000",56994 => "0000000000000000",
56995 => "0000000000000000",56996 => "0000000000000000",
56997 => "0000000000000000",56998 => "0000000000000000",
56999 => "0000000000000000",57000 => "0000000000000000",
57001 => "0000000000000000",57002 => "0000000000000000",
57003 => "0000000000000000",57004 => "0000000000000000",
57005 => "0000000000000000",57006 => "0000000000000000",
57007 => "0000000000000000",57008 => "0000000000000000",
57009 => "0000000000000000",57010 => "0000000000000000",
57011 => "0000000000000000",57012 => "0000000000000000",
57013 => "0000000000000000",57014 => "0000000000000000",
57015 => "0000000000000000",57016 => "0000000000000000",
57017 => "0000000000000000",57018 => "0000000000000000",
57019 => "0000000000000000",57020 => "0000000000000000",
57021 => "0000000000000000",57022 => "0000000000000000",
57023 => "0000000000000000",57024 => "0000000000000000",
57025 => "0000000000000000",57026 => "0000000000000000",
57027 => "0000000000000000",57028 => "0000000000000000",
57029 => "0000000000000000",57030 => "0000000000000000",
57031 => "0000000000000000",57032 => "0000000000000000",
57033 => "0000000000000000",57034 => "0000000000000000",
57035 => "0000000000000000",57036 => "0000000000000000",
57037 => "0000000000000000",57038 => "0000000000000000",
57039 => "0000000000000000",57040 => "0000000000000000",
57041 => "0000000000000000",57042 => "0000000000000000",
57043 => "0000000000000000",57044 => "0000000000000000",
57045 => "0000000000000000",57046 => "0000000000000000",
57047 => "0000000000000000",57048 => "0000000000000000",
57049 => "0000000000000000",57050 => "0000000000000000",
57051 => "0000000000000000",57052 => "0000000000000000",
57053 => "0000000000000000",57054 => "0000000000000000",
57055 => "0000000000000000",57056 => "0000000000000000",
57057 => "0000000000000000",57058 => "0000000000000000",
57059 => "0000000000000000",57060 => "0000000000000000",
57061 => "0000000000000000",57062 => "0000000000000000",
57063 => "0000000000000000",57064 => "0000000000000000",
57065 => "0000000000000000",57066 => "0000000000000000",
57067 => "0000000000000000",57068 => "0000000000000000",
57069 => "0000000000000000",57070 => "0000000000000000",
57071 => "0000000000000000",57072 => "0000000000000000",
57073 => "0000000000000000",57074 => "0000000000000000",
57075 => "0000000000000000",57076 => "0000000000000000",
57077 => "0000000000000000",57078 => "0000000000000000",
57079 => "0000000000000000",57080 => "0000000000000000",
57081 => "0000000000000000",57082 => "0000000000000000",
57083 => "0000000000000000",57084 => "0000000000000000",
57085 => "0000000000000000",57086 => "0000000000000000",
57087 => "0000000000000000",57088 => "0000000000000000",
57089 => "0000000000000000",57090 => "0000000000000000",
57091 => "0000000000000000",57092 => "0000000000000000",
57093 => "0000000000000000",57094 => "0000000000000000",
57095 => "0000000000000000",57096 => "0000000000000000",
57097 => "0000000000000000",57098 => "0000000000000000",
57099 => "0000000000000000",57100 => "0000000000000000",
57101 => "0000000000000000",57102 => "0000000000000000",
57103 => "0000000000000000",57104 => "0000000000000000",
57105 => "0000000000000000",57106 => "0000000000000000",
57107 => "0000000000000000",57108 => "0000000000000000",
57109 => "0000000000000000",57110 => "0000000000000000",
57111 => "0000000000000000",57112 => "0000000000000000",
57113 => "0000000000000000",57114 => "0000000000000000",
57115 => "0000000000000000",57116 => "0000000000000000",
57117 => "0000000000000000",57118 => "0000000000000000",
57119 => "0000000000000000",57120 => "0000000000000000",
57121 => "0000000000000000",57122 => "0000000000000000",
57123 => "0000000000000000",57124 => "0000000000000000",
57125 => "0000000000000000",57126 => "0000000000000000",
57127 => "0000000000000000",57128 => "0000000000000000",
57129 => "0000000000000000",57130 => "0000000000000000",
57131 => "0000000000000000",57132 => "0000000000000000",
57133 => "0000000000000000",57134 => "0000000000000000",
57135 => "0000000000000000",57136 => "0000000000000000",
57137 => "0000000000000000",57138 => "0000000000000000",
57139 => "0000000000000000",57140 => "0000000000000000",
57141 => "0000000000000000",57142 => "0000000000000000",
57143 => "0000000000000000",57144 => "0000000000000000",
57145 => "0000000000000000",57146 => "0000000000000000",
57147 => "0000000000000000",57148 => "0000000000000000",
57149 => "0000000000000000",57150 => "0000000000000000",
57151 => "0000000000000000",57152 => "0000000000000000",
57153 => "0000000000000000",57154 => "0000000000000000",
57155 => "0000000000000000",57156 => "0000000000000000",
57157 => "0000000000000000",57158 => "0000000000000000",
57159 => "0000000000000000",57160 => "0000000000000000",
57161 => "0000000000000000",57162 => "0000000000000000",
57163 => "0000000000000000",57164 => "0000000000000000",
57165 => "0000000000000000",57166 => "0000000000000000",
57167 => "0000000000000000",57168 => "0000000000000000",
57169 => "0000000000000000",57170 => "0000000000000000",
57171 => "0000000000000000",57172 => "0000000000000000",
57173 => "0000000000000000",57174 => "0000000000000000",
57175 => "0000000000000000",57176 => "0000000000000000",
57177 => "0000000000000000",57178 => "0000000000000000",
57179 => "0000000000000000",57180 => "0000000000000000",
57181 => "0000000000000000",57182 => "0000000000000000",
57183 => "0000000000000000",57184 => "0000000000000000",
57185 => "0000000000000000",57186 => "0000000000000000",
57187 => "0000000000000000",57188 => "0000000000000000",
57189 => "0000000000000000",57190 => "0000000000000000",
57191 => "0000000000000000",57192 => "0000000000000000",
57193 => "0000000000000000",57194 => "0000000000000000",
57195 => "0000000000000000",57196 => "0000000000000000",
57197 => "0000000000000000",57198 => "0000000000000000",
57199 => "0000000000000000",57200 => "0000000000000000",
57201 => "0000000000000000",57202 => "0000000000000000",
57203 => "0000000000000000",57204 => "0000000000000000",
57205 => "0000000000000000",57206 => "0000000000000000",
57207 => "0000000000000000",57208 => "0000000000000000",
57209 => "0000000000000000",57210 => "0000000000000000",
57211 => "0000000000000000",57212 => "0000000000000000",
57213 => "0000000000000000",57214 => "0000000000000000",
57215 => "0000000000000000",57216 => "0000000000000000",
57217 => "0000000000000000",57218 => "0000000000000000",
57219 => "0000000000000000",57220 => "0000000000000000",
57221 => "0000000000000000",57222 => "0000000000000000",
57223 => "0000000000000000",57224 => "0000000000000000",
57225 => "0000000000000000",57226 => "0000000000000000",
57227 => "0000000000000000",57228 => "0000000000000000",
57229 => "0000000000000000",57230 => "0000000000000000",
57231 => "0000000000000000",57232 => "0000000000000000",
57233 => "0000000000000000",57234 => "0000000000000000",
57235 => "0000000000000000",57236 => "0000000000000000",
57237 => "0000000000000000",57238 => "0000000000000000",
57239 => "0000000000000000",57240 => "0000000000000000",
57241 => "0000000000000000",57242 => "0000000000000000",
57243 => "0000000000000000",57244 => "0000000000000000",
57245 => "0000000000000000",57246 => "0000000000000000",
57247 => "0000000000000000",57248 => "0000000000000000",
57249 => "0000000000000000",57250 => "0000000000000000",
57251 => "0000000000000000",57252 => "0000000000000000",
57253 => "0000000000000000",57254 => "0000000000000000",
57255 => "0000000000000000",57256 => "0000000000000000",
57257 => "0000000000000000",57258 => "0000000000000000",
57259 => "0000000000000000",57260 => "0000000000000000",
57261 => "0000000000000000",57262 => "0000000000000000",
57263 => "0000000000000000",57264 => "0000000000000000",
57265 => "0000000000000000",57266 => "0000000000000000",
57267 => "0000000000000000",57268 => "0000000000000000",
57269 => "0000000000000000",57270 => "0000000000000000",
57271 => "0000000000000000",57272 => "0000000000000000",
57273 => "0000000000000000",57274 => "0000000000000000",
57275 => "0000000000000000",57276 => "0000000000000000",
57277 => "0000000000000000",57278 => "0000000000000000",
57279 => "0000000000000000",57280 => "0000000000000000",
57281 => "0000000000000000",57282 => "0000000000000000",
57283 => "0000000000000000",57284 => "0000000000000000",
57285 => "0000000000000000",57286 => "0000000000000000",
57287 => "0000000000000000",57288 => "0000000000000000",
57289 => "0000000000000000",57290 => "0000000000000000",
57291 => "0000000000000000",57292 => "0000000000000000",
57293 => "0000000000000000",57294 => "0000000000000000",
57295 => "0000000000000000",57296 => "0000000000000000",
57297 => "0000000000000000",57298 => "0000000000000000",
57299 => "0000000000000000",57300 => "0000000000000000",
57301 => "0000000000000000",57302 => "0000000000000000",
57303 => "0000000000000000",57304 => "0000000000000000",
57305 => "0000000000000000",57306 => "0000000000000000",
57307 => "0000000000000000",57308 => "0000000000000000",
57309 => "0000000000000000",57310 => "0000000000000000",
57311 => "0000000000000000",57312 => "0000000000000000",
57313 => "0000000000000000",57314 => "0000000000000000",
57315 => "0000000000000000",57316 => "0000000000000000",
57317 => "0000000000000000",57318 => "0000000000000000",
57319 => "0000000000000000",57320 => "0000000000000000",
57321 => "0000000000000000",57322 => "0000000000000000",
57323 => "0000000000000000",57324 => "0000000000000000",
57325 => "0000000000000000",57326 => "0000000000000000",
57327 => "0000000000000000",57328 => "0000000000000000",
57329 => "0000000000000000",57330 => "0000000000000000",
57331 => "0000000000000000",57332 => "0000000000000000",
57333 => "0000000000000000",57334 => "0000000000000000",
57335 => "0000000000000000",57336 => "0000000000000000",
57337 => "0000000000000000",57338 => "0000000000000000",
57339 => "0000000000000000",57340 => "0000000000000000",
57341 => "0000000000000000",57342 => "0000000000000000",
57343 => "0000000000000000",57344 => "0000000000000000",
57345 => "0000000000000000",57346 => "0000000000000000",
57347 => "0000000000000000",57348 => "0000000000000000",
57349 => "0000000000000000",57350 => "0000000000000000",
57351 => "0000000000000000",57352 => "0000000000000000",
57353 => "0000000000000000",57354 => "0000000000000000",
57355 => "0000000000000000",57356 => "0000000000000000",
57357 => "0000000000000000",57358 => "0000000000000000",
57359 => "0000000000000000",57360 => "0000000000000000",
57361 => "0000000000000000",57362 => "0000000000000000",
57363 => "0000000000000000",57364 => "0000000000000000",
57365 => "0000000000000000",57366 => "0000000000000000",
57367 => "0000000000000000",57368 => "0000000000000000",
57369 => "0000000000000000",57370 => "0000000000000000",
57371 => "0000000000000000",57372 => "0000000000000000",
57373 => "0000000000000000",57374 => "0000000000000000",
57375 => "0000000000000000",57376 => "0000000000000000",
57377 => "0000000000000000",57378 => "0000000000000000",
57379 => "0000000000000000",57380 => "0000000000000000",
57381 => "0000000000000000",57382 => "0000000000000000",
57383 => "0000000000000000",57384 => "0000000000000000",
57385 => "0000000000000000",57386 => "0000000000000000",
57387 => "0000000000000000",57388 => "0000000000000000",
57389 => "0000000000000000",57390 => "0000000000000000",
57391 => "0000000000000000",57392 => "0000000000000000",
57393 => "0000000000000000",57394 => "0000000000000000",
57395 => "0000000000000000",57396 => "0000000000000000",
57397 => "0000000000000000",57398 => "0000000000000000",
57399 => "0000000000000000",57400 => "0000000000000000",
57401 => "0000000000000000",57402 => "0000000000000000",
57403 => "0000000000000000",57404 => "0000000000000000",
57405 => "0000000000000000",57406 => "0000000000000000",
57407 => "0000000000000000",57408 => "0000000000000000",
57409 => "0000000000000000",57410 => "0000000000000000",
57411 => "0000000000000000",57412 => "0000000000000000",
57413 => "0000000000000000",57414 => "0000000000000000",
57415 => "0000000000000000",57416 => "0000000000000000",
57417 => "0000000000000000",57418 => "0000000000000000",
57419 => "0000000000000000",57420 => "0000000000000000",
57421 => "0000000000000000",57422 => "0000000000000000",
57423 => "0000000000000000",57424 => "0000000000000000",
57425 => "0000000000000000",57426 => "0000000000000000",
57427 => "0000000000000000",57428 => "0000000000000000",
57429 => "0000000000000000",57430 => "0000000000000000",
57431 => "0000000000000000",57432 => "0000000000000000",
57433 => "0000000000000000",57434 => "0000000000000000",
57435 => "0000000000000000",57436 => "0000000000000000",
57437 => "0000000000000000",57438 => "0000000000000000",
57439 => "0000000000000000",57440 => "0000000000000000",
57441 => "0000000000000000",57442 => "0000000000000000",
57443 => "0000000000000000",57444 => "0000000000000000",
57445 => "0000000000000000",57446 => "0000000000000000",
57447 => "0000000000000000",57448 => "0000000000000000",
57449 => "0000000000000000",57450 => "0000000000000000",
57451 => "0000000000000000",57452 => "0000000000000000",
57453 => "0000000000000000",57454 => "0000000000000000",
57455 => "0000000000000000",57456 => "0000000000000000",
57457 => "0000000000000000",57458 => "0000000000000000",
57459 => "0000000000000000",57460 => "0000000000000000",
57461 => "0000000000000000",57462 => "0000000000000000",
57463 => "0000000000000000",57464 => "0000000000000000",
57465 => "0000000000000000",57466 => "0000000000000000",
57467 => "0000000000000000",57468 => "0000000000000000",
57469 => "0000000000000000",57470 => "0000000000000000",
57471 => "0000000000000000",57472 => "0000000000000000",
57473 => "0000000000000000",57474 => "0000000000000000",
57475 => "0000000000000000",57476 => "0000000000000000",
57477 => "0000000000000000",57478 => "0000000000000000",
57479 => "0000000000000000",57480 => "0000000000000000",
57481 => "0000000000000000",57482 => "0000000000000000",
57483 => "0000000000000000",57484 => "0000000000000000",
57485 => "0000000000000000",57486 => "0000000000000000",
57487 => "0000000000000000",57488 => "0000000000000000",
57489 => "0000000000000000",57490 => "0000000000000000",
57491 => "0000000000000000",57492 => "0000000000000000",
57493 => "0000000000000000",57494 => "0000000000000000",
57495 => "0000000000000000",57496 => "0000000000000000",
57497 => "0000000000000000",57498 => "0000000000000000",
57499 => "0000000000000000",57500 => "0000000000000000",
57501 => "0000000000000000",57502 => "0000000000000000",
57503 => "0000000000000000",57504 => "0000000000000000",
57505 => "0000000000000000",57506 => "0000000000000000",
57507 => "0000000000000000",57508 => "0000000000000000",
57509 => "0000000000000000",57510 => "0000000000000000",
57511 => "0000000000000000",57512 => "0000000000000000",
57513 => "0000000000000000",57514 => "0000000000000000",
57515 => "0000000000000000",57516 => "0000000000000000",
57517 => "0000000000000000",57518 => "0000000000000000",
57519 => "0000000000000000",57520 => "0000000000000000",
57521 => "0000000000000000",57522 => "0000000000000000",
57523 => "0000000000000000",57524 => "0000000000000000",
57525 => "0000000000000000",57526 => "0000000000000000",
57527 => "0000000000000000",57528 => "0000000000000000",
57529 => "0000000000000000",57530 => "0000000000000000",
57531 => "0000000000000000",57532 => "0000000000000000",
57533 => "0000000000000000",57534 => "0000000000000000",
57535 => "0000000000000000",57536 => "0000000000000000",
57537 => "0000000000000000",57538 => "0000000000000000",
57539 => "0000000000000000",57540 => "0000000000000000",
57541 => "0000000000000000",57542 => "0000000000000000",
57543 => "0000000000000000",57544 => "0000000000000000",
57545 => "0000000000000000",57546 => "0000000000000000",
57547 => "0000000000000000",57548 => "0000000000000000",
57549 => "0000000000000000",57550 => "0000000000000000",
57551 => "0000000000000000",57552 => "0000000000000000",
57553 => "0000000000000000",57554 => "0000000000000000",
57555 => "0000000000000000",57556 => "0000000000000000",
57557 => "0000000000000000",57558 => "0000000000000000",
57559 => "0000000000000000",57560 => "0000000000000000",
57561 => "0000000000000000",57562 => "0000000000000000",
57563 => "0000000000000000",57564 => "0000000000000000",
57565 => "0000000000000000",57566 => "0000000000000000",
57567 => "0000000000000000",57568 => "0000000000000000",
57569 => "0000000000000000",57570 => "0000000000000000",
57571 => "0000000000000000",57572 => "0000000000000000",
57573 => "0000000000000000",57574 => "0000000000000000",
57575 => "0000000000000000",57576 => "0000000000000000",
57577 => "0000000000000000",57578 => "0000000000000000",
57579 => "0000000000000000",57580 => "0000000000000000",
57581 => "0000000000000000",57582 => "0000000000000000",
57583 => "0000000000000000",57584 => "0000000000000000",
57585 => "0000000000000000",57586 => "0000000000000000",
57587 => "0000000000000000",57588 => "0000000000000000",
57589 => "0000000000000000",57590 => "0000000000000000",
57591 => "0000000000000000",57592 => "0000000000000000",
57593 => "0000000000000000",57594 => "0000000000000000",
57595 => "0000000000000000",57596 => "0000000000000000",
57597 => "0000000000000000",57598 => "0000000000000000",
57599 => "0000000000000000",57600 => "0000000000000000",
57601 => "0000000000000000",57602 => "0000000000000000",
57603 => "0000000000000000",57604 => "0000000000000000",
57605 => "0000000000000000",57606 => "0000000000000000",
57607 => "0000000000000000",57608 => "0000000000000000",
57609 => "0000000000000000",57610 => "0000000000000000",
57611 => "0000000000000000",57612 => "0000000000000000",
57613 => "0000000000000000",57614 => "0000000000000000",
57615 => "0000000000000000",57616 => "0000000000000000",
57617 => "0000000000000000",57618 => "0000000000000000",
57619 => "0000000000000000",57620 => "0000000000000000",
57621 => "0000000000000000",57622 => "0000000000000000",
57623 => "0000000000000000",57624 => "0000000000000000",
57625 => "0000000000000000",57626 => "0000000000000000",
57627 => "0000000000000000",57628 => "0000000000000000",
57629 => "0000000000000000",57630 => "0000000000000000",
57631 => "0000000000000000",57632 => "0000000000000000",
57633 => "0000000000000000",57634 => "0000000000000000",
57635 => "0000000000000000",57636 => "0000000000000000",
57637 => "0000000000000000",57638 => "0000000000000000",
57639 => "0000000000000000",57640 => "0000000000000000",
57641 => "0000000000000000",57642 => "0000000000000000",
57643 => "0000000000000000",57644 => "0000000000000000",
57645 => "0000000000000000",57646 => "0000000000000000",
57647 => "0000000000000000",57648 => "0000000000000000",
57649 => "0000000000000000",57650 => "0000000000000000",
57651 => "0000000000000000",57652 => "0000000000000000",
57653 => "0000000000000000",57654 => "0000000000000000",
57655 => "0000000000000000",57656 => "0000000000000000",
57657 => "0000000000000000",57658 => "0000000000000000",
57659 => "0000000000000000",57660 => "0000000000000000",
57661 => "0000000000000000",57662 => "0000000000000000",
57663 => "0000000000000000",57664 => "0000000000000000",
57665 => "0000000000000000",57666 => "0000000000000000",
57667 => "0000000000000000",57668 => "0000000000000000",
57669 => "0000000000000000",57670 => "0000000000000000",
57671 => "0000000000000000",57672 => "0000000000000000",
57673 => "0000000000000000",57674 => "0000000000000000",
57675 => "0000000000000000",57676 => "0000000000000000",
57677 => "0000000000000000",57678 => "0000000000000000",
57679 => "0000000000000000",57680 => "0000000000000000",
57681 => "0000000000000000",57682 => "0000000000000000",
57683 => "0000000000000000",57684 => "0000000000000000",
57685 => "0000000000000000",57686 => "0000000000000000",
57687 => "0000000000000000",57688 => "0000000000000000",
57689 => "0000000000000000",57690 => "0000000000000000",
57691 => "0000000000000000",57692 => "0000000000000000",
57693 => "0000000000000000",57694 => "0000000000000000",
57695 => "0000000000000000",57696 => "0000000000000000",
57697 => "0000000000000000",57698 => "0000000000000000",
57699 => "0000000000000000",57700 => "0000000000000000",
57701 => "0000000000000000",57702 => "0000000000000000",
57703 => "0000000000000000",57704 => "0000000000000000",
57705 => "0000000000000000",57706 => "0000000000000000",
57707 => "0000000000000000",57708 => "0000000000000000",
57709 => "0000000000000000",57710 => "0000000000000000",
57711 => "0000000000000000",57712 => "0000000000000000",
57713 => "0000000000000000",57714 => "0000000000000000",
57715 => "0000000000000000",57716 => "0000000000000000",
57717 => "0000000000000000",57718 => "0000000000000000",
57719 => "0000000000000000",57720 => "0000000000000000",
57721 => "0000000000000000",57722 => "0000000000000000",
57723 => "0000000000000000",57724 => "0000000000000000",
57725 => "0000000000000000",57726 => "0000000000000000",
57727 => "0000000000000000",57728 => "0000000000000000",
57729 => "0000000000000000",57730 => "0000000000000000",
57731 => "0000000000000000",57732 => "0000000000000000",
57733 => "0000000000000000",57734 => "0000000000000000",
57735 => "0000000000000000",57736 => "0000000000000000",
57737 => "0000000000000000",57738 => "0000000000000000",
57739 => "0000000000000000",57740 => "0000000000000000",
57741 => "0000000000000000",57742 => "0000000000000000",
57743 => "0000000000000000",57744 => "0000000000000000",
57745 => "0000000000000000",57746 => "0000000000000000",
57747 => "0000000000000000",57748 => "0000000000000000",
57749 => "0000000000000000",57750 => "0000000000000000",
57751 => "0000000000000000",57752 => "0000000000000000",
57753 => "0000000000000000",57754 => "0000000000000000",
57755 => "0000000000000000",57756 => "0000000000000000",
57757 => "0000000000000000",57758 => "0000000000000000",
57759 => "0000000000000000",57760 => "0000000000000000",
57761 => "0000000000000000",57762 => "0000000000000000",
57763 => "0000000000000000",57764 => "0000000000000000",
57765 => "0000000000000000",57766 => "0000000000000000",
57767 => "0000000000000000",57768 => "0000000000000000",
57769 => "0000000000000000",57770 => "0000000000000000",
57771 => "0000000000000000",57772 => "0000000000000000",
57773 => "0000000000000000",57774 => "0000000000000000",
57775 => "0000000000000000",57776 => "0000000000000000",
57777 => "0000000000000000",57778 => "0000000000000000",
57779 => "0000000000000000",57780 => "0000000000000000",
57781 => "0000000000000000",57782 => "0000000000000000",
57783 => "0000000000000000",57784 => "0000000000000000",
57785 => "0000000000000000",57786 => "0000000000000000",
57787 => "0000000000000000",57788 => "0000000000000000",
57789 => "0000000000000000",57790 => "0000000000000000",
57791 => "0000000000000000",57792 => "0000000000000000",
57793 => "0000000000000000",57794 => "0000000000000000",
57795 => "0000000000000000",57796 => "0000000000000000",
57797 => "0000000000000000",57798 => "0000000000000000",
57799 => "0000000000000000",57800 => "0000000000000000",
57801 => "0000000000000000",57802 => "0000000000000000",
57803 => "0000000000000000",57804 => "0000000000000000",
57805 => "0000000000000000",57806 => "0000000000000000",
57807 => "0000000000000000",57808 => "0000000000000000",
57809 => "0000000000000000",57810 => "0000000000000000",
57811 => "0000000000000000",57812 => "0000000000000000",
57813 => "0000000000000000",57814 => "0000000000000000",
57815 => "0000000000000000",57816 => "0000000000000000",
57817 => "0000000000000000",57818 => "0000000000000000",
57819 => "0000000000000000",57820 => "0000000000000000",
57821 => "0000000000000000",57822 => "0000000000000000",
57823 => "0000000000000000",57824 => "0000000000000000",
57825 => "0000000000000000",57826 => "0000000000000000",
57827 => "0000000000000000",57828 => "0000000000000000",
57829 => "0000000000000000",57830 => "0000000000000000",
57831 => "0000000000000000",57832 => "0000000000000000",
57833 => "0000000000000000",57834 => "0000000000000000",
57835 => "0000000000000000",57836 => "0000000000000000",
57837 => "0000000000000000",57838 => "0000000000000000",
57839 => "0000000000000000",57840 => "0000000000000000",
57841 => "0000000000000000",57842 => "0000000000000000",
57843 => "0000000000000000",57844 => "0000000000000000",
57845 => "0000000000000000",57846 => "0000000000000000",
57847 => "0000000000000000",57848 => "0000000000000000",
57849 => "0000000000000000",57850 => "0000000000000000",
57851 => "0000000000000000",57852 => "0000000000000000",
57853 => "0000000000000000",57854 => "0000000000000000",
57855 => "0000000000000000",57856 => "0000000000000000",
57857 => "0000000000000000",57858 => "0000000000000000",
57859 => "0000000000000000",57860 => "0000000000000000",
57861 => "0000000000000000",57862 => "0000000000000000",
57863 => "0000000000000000",57864 => "0000000000000000",
57865 => "0000000000000000",57866 => "0000000000000000",
57867 => "0000000000000000",57868 => "0000000000000000",
57869 => "0000000000000000",57870 => "0000000000000000",
57871 => "0000000000000000",57872 => "0000000000000000",
57873 => "0000000000000000",57874 => "0000000000000000",
57875 => "0000000000000000",57876 => "0000000000000000",
57877 => "0000000000000000",57878 => "0000000000000000",
57879 => "0000000000000000",57880 => "0000000000000000",
57881 => "0000000000000000",57882 => "0000000000000000",
57883 => "0000000000000000",57884 => "0000000000000000",
57885 => "0000000000000000",57886 => "0000000000000000",
57887 => "0000000000000000",57888 => "0000000000000000",
57889 => "0000000000000000",57890 => "0000000000000000",
57891 => "0000000000000000",57892 => "0000000000000000",
57893 => "0000000000000000",57894 => "0000000000000000",
57895 => "0000000000000000",57896 => "0000000000000000",
57897 => "0000000000000000",57898 => "0000000000000000",
57899 => "0000000000000000",57900 => "0000000000000000",
57901 => "0000000000000000",57902 => "0000000000000000",
57903 => "0000000000000000",57904 => "0000000000000000",
57905 => "0000000000000000",57906 => "0000000000000000",
57907 => "0000000000000000",57908 => "0000000000000000",
57909 => "0000000000000000",57910 => "0000000000000000",
57911 => "0000000000000000",57912 => "0000000000000000",
57913 => "0000000000000000",57914 => "0000000000000000",
57915 => "0000000000000000",57916 => "0000000000000000",
57917 => "0000000000000000",57918 => "0000000000000000",
57919 => "0000000000000000",57920 => "0000000000000000",
57921 => "0000000000000000",57922 => "0000000000000000",
57923 => "0000000000000000",57924 => "0000000000000000",
57925 => "0000000000000000",57926 => "0000000000000000",
57927 => "0000000000000000",57928 => "0000000000000000",
57929 => "0000000000000000",57930 => "0000000000000000",
57931 => "0000000000000000",57932 => "0000000000000000",
57933 => "0000000000000000",57934 => "0000000000000000",
57935 => "0000000000000000",57936 => "0000000000000000",
57937 => "0000000000000000",57938 => "0000000000000000",
57939 => "0000000000000000",57940 => "0000000000000000",
57941 => "0000000000000000",57942 => "0000000000000000",
57943 => "0000000000000000",57944 => "0000000000000000",
57945 => "0000000000000000",57946 => "0000000000000000",
57947 => "0000000000000000",57948 => "0000000000000000",
57949 => "0000000000000000",57950 => "0000000000000000",
57951 => "0000000000000000",57952 => "0000000000000000",
57953 => "0000000000000000",57954 => "0000000000000000",
57955 => "0000000000000000",57956 => "0000000000000000",
57957 => "0000000000000000",57958 => "0000000000000000",
57959 => "0000000000000000",57960 => "0000000000000000",
57961 => "0000000000000000",57962 => "0000000000000000",
57963 => "0000000000000000",57964 => "0000000000000000",
57965 => "0000000000000000",57966 => "0000000000000000",
57967 => "0000000000000000",57968 => "0000000000000000",
57969 => "0000000000000000",57970 => "0000000000000000",
57971 => "0000000000000000",57972 => "0000000000000000",
57973 => "0000000000000000",57974 => "0000000000000000",
57975 => "0000000000000000",57976 => "0000000000000000",
57977 => "0000000000000000",57978 => "0000000000000000",
57979 => "0000000000000000",57980 => "0000000000000000",
57981 => "0000000000000000",57982 => "0000000000000000",
57983 => "0000000000000000",57984 => "0000000000000000",
57985 => "0000000000000000",57986 => "0000000000000000",
57987 => "0000000000000000",57988 => "0000000000000000",
57989 => "0000000000000000",57990 => "0000000000000000",
57991 => "0000000000000000",57992 => "0000000000000000",
57993 => "0000000000000000",57994 => "0000000000000000",
57995 => "0000000000000000",57996 => "0000000000000000",
57997 => "0000000000000000",57998 => "0000000000000000",
57999 => "0000000000000000",58000 => "0000000000000000",
58001 => "0000000000000000",58002 => "0000000000000000",
58003 => "0000000000000000",58004 => "0000000000000000",
58005 => "0000000000000000",58006 => "0000000000000000",
58007 => "0000000000000000",58008 => "0000000000000000",
58009 => "0000000000000000",58010 => "0000000000000000",
58011 => "0000000000000000",58012 => "0000000000000000",
58013 => "0000000000000000",58014 => "0000000000000000",
58015 => "0000000000000000",58016 => "0000000000000000",
58017 => "0000000000000000",58018 => "0000000000000000",
58019 => "0000000000000000",58020 => "0000000000000000",
58021 => "0000000000000000",58022 => "0000000000000000",
58023 => "0000000000000000",58024 => "0000000000000000",
58025 => "0000000000000000",58026 => "0000000000000000",
58027 => "0000000000000000",58028 => "0000000000000000",
58029 => "0000000000000000",58030 => "0000000000000000",
58031 => "0000000000000000",58032 => "0000000000000000",
58033 => "0000000000000000",58034 => "0000000000000000",
58035 => "0000000000000000",58036 => "0000000000000000",
58037 => "0000000000000000",58038 => "0000000000000000",
58039 => "0000000000000000",58040 => "0000000000000000",
58041 => "0000000000000000",58042 => "0000000000000000",
58043 => "0000000000000000",58044 => "0000000000000000",
58045 => "0000000000000000",58046 => "0000000000000000",
58047 => "0000000000000000",58048 => "0000000000000000",
58049 => "0000000000000000",58050 => "0000000000000000",
58051 => "0000000000000000",58052 => "0000000000000000",
58053 => "0000000000000000",58054 => "0000000000000000",
58055 => "0000000000000000",58056 => "0000000000000000",
58057 => "0000000000000000",58058 => "0000000000000000",
58059 => "0000000000000000",58060 => "0000000000000000",
58061 => "0000000000000000",58062 => "0000000000000000",
58063 => "0000000000000000",58064 => "0000000000000000",
58065 => "0000000000000000",58066 => "0000000000000000",
58067 => "0000000000000000",58068 => "0000000000000000",
58069 => "0000000000000000",58070 => "0000000000000000",
58071 => "0000000000000000",58072 => "0000000000000000",
58073 => "0000000000000000",58074 => "0000000000000000",
58075 => "0000000000000000",58076 => "0000000000000000",
58077 => "0000000000000000",58078 => "0000000000000000",
58079 => "0000000000000000",58080 => "0000000000000000",
58081 => "0000000000000000",58082 => "0000000000000000",
58083 => "0000000000000000",58084 => "0000000000000000",
58085 => "0000000000000000",58086 => "0000000000000000",
58087 => "0000000000000000",58088 => "0000000000000000",
58089 => "0000000000000000",58090 => "0000000000000000",
58091 => "0000000000000000",58092 => "0000000000000000",
58093 => "0000000000000000",58094 => "0000000000000000",
58095 => "0000000000000000",58096 => "0000000000000000",
58097 => "0000000000000000",58098 => "0000000000000000",
58099 => "0000000000000000",58100 => "0000000000000000",
58101 => "0000000000000000",58102 => "0000000000000000",
58103 => "0000000000000000",58104 => "0000000000000000",
58105 => "0000000000000000",58106 => "0000000000000000",
58107 => "0000000000000000",58108 => "0000000000000000",
58109 => "0000000000000000",58110 => "0000000000000000",
58111 => "0000000000000000",58112 => "0000000000000000",
58113 => "0000000000000000",58114 => "0000000000000000",
58115 => "0000000000000000",58116 => "0000000000000000",
58117 => "0000000000000000",58118 => "0000000000000000",
58119 => "0000000000000000",58120 => "0000000000000000",
58121 => "0000000000000000",58122 => "0000000000000000",
58123 => "0000000000000000",58124 => "0000000000000000",
58125 => "0000000000000000",58126 => "0000000000000000",
58127 => "0000000000000000",58128 => "0000000000000000",
58129 => "0000000000000000",58130 => "0000000000000000",
58131 => "0000000000000000",58132 => "0000000000000000",
58133 => "0000000000000000",58134 => "0000000000000000",
58135 => "0000000000000000",58136 => "0000000000000000",
58137 => "0000000000000000",58138 => "0000000000000000",
58139 => "0000000000000000",58140 => "0000000000000000",
58141 => "0000000000000000",58142 => "0000000000000000",
58143 => "0000000000000000",58144 => "0000000000000000",
58145 => "0000000000000000",58146 => "0000000000000000",
58147 => "0000000000000000",58148 => "0000000000000000",
58149 => "0000000000000000",58150 => "0000000000000000",
58151 => "0000000000000000",58152 => "0000000000000000",
58153 => "0000000000000000",58154 => "0000000000000000",
58155 => "0000000000000000",58156 => "0000000000000000",
58157 => "0000000000000000",58158 => "0000000000000000",
58159 => "0000000000000000",58160 => "0000000000000000",
58161 => "0000000000000000",58162 => "0000000000000000",
58163 => "0000000000000000",58164 => "0000000000000000",
58165 => "0000000000000000",58166 => "0000000000000000",
58167 => "0000000000000000",58168 => "0000000000000000",
58169 => "0000000000000000",58170 => "0000000000000000",
58171 => "0000000000000000",58172 => "0000000000000000",
58173 => "0000000000000000",58174 => "0000000000000000",
58175 => "0000000000000000",58176 => "0000000000000000",
58177 => "0000000000000000",58178 => "0000000000000000",
58179 => "0000000000000000",58180 => "0000000000000000",
58181 => "0000000000000000",58182 => "0000000000000000",
58183 => "0000000000000000",58184 => "0000000000000000",
58185 => "0000000000000000",58186 => "0000000000000000",
58187 => "0000000000000000",58188 => "0000000000000000",
58189 => "0000000000000000",58190 => "0000000000000000",
58191 => "0000000000000000",58192 => "0000000000000000",
58193 => "0000000000000000",58194 => "0000000000000000",
58195 => "0000000000000000",58196 => "0000000000000000",
58197 => "0000000000000000",58198 => "0000000000000000",
58199 => "0000000000000000",58200 => "0000000000000000",
58201 => "0000000000000000",58202 => "0000000000000000",
58203 => "0000000000000000",58204 => "0000000000000000",
58205 => "0000000000000000",58206 => "0000000000000000",
58207 => "0000000000000000",58208 => "0000000000000000",
58209 => "0000000000000000",58210 => "0000000000000000",
58211 => "0000000000000000",58212 => "0000000000000000",
58213 => "0000000000000000",58214 => "0000000000000000",
58215 => "0000000000000000",58216 => "0000000000000000",
58217 => "0000000000000000",58218 => "0000000000000000",
58219 => "0000000000000000",58220 => "0000000000000000",
58221 => "0000000000000000",58222 => "0000000000000000",
58223 => "0000000000000000",58224 => "0000000000000000",
58225 => "0000000000000000",58226 => "0000000000000000",
58227 => "0000000000000000",58228 => "0000000000000000",
58229 => "0000000000000000",58230 => "0000000000000000",
58231 => "0000000000000000",58232 => "0000000000000000",
58233 => "0000000000000000",58234 => "0000000000000000",
58235 => "0000000000000000",58236 => "0000000000000000",
58237 => "0000000000000000",58238 => "0000000000000000",
58239 => "0000000000000000",58240 => "0000000000000000",
58241 => "0000000000000000",58242 => "0000000000000000",
58243 => "0000000000000000",58244 => "0000000000000000",
58245 => "0000000000000000",58246 => "0000000000000000",
58247 => "0000000000000000",58248 => "0000000000000000",
58249 => "0000000000000000",58250 => "0000000000000000",
58251 => "0000000000000000",58252 => "0000000000000000",
58253 => "0000000000000000",58254 => "0000000000000000",
58255 => "0000000000000000",58256 => "0000000000000000",
58257 => "0000000000000000",58258 => "0000000000000000",
58259 => "0000000000000000",58260 => "0000000000000000",
58261 => "0000000000000000",58262 => "0000000000000000",
58263 => "0000000000000000",58264 => "0000000000000000",
58265 => "0000000000000000",58266 => "0000000000000000",
58267 => "0000000000000000",58268 => "0000000000000000",
58269 => "0000000000000000",58270 => "0000000000000000",
58271 => "0000000000000000",58272 => "0000000000000000",
58273 => "0000000000000000",58274 => "0000000000000000",
58275 => "0000000000000000",58276 => "0000000000000000",
58277 => "0000000000000000",58278 => "0000000000000000",
58279 => "0000000000000000",58280 => "0000000000000000",
58281 => "0000000000000000",58282 => "0000000000000000",
58283 => "0000000000000000",58284 => "0000000000000000",
58285 => "0000000000000000",58286 => "0000000000000000",
58287 => "0000000000000000",58288 => "0000000000000000",
58289 => "0000000000000000",58290 => "0000000000000000",
58291 => "0000000000000000",58292 => "0000000000000000",
58293 => "0000000000000000",58294 => "0000000000000000",
58295 => "0000000000000000",58296 => "0000000000000000",
58297 => "0000000000000000",58298 => "0000000000000000",
58299 => "0000000000000000",58300 => "0000000000000000",
58301 => "0000000000000000",58302 => "0000000000000000",
58303 => "0000000000000000",58304 => "0000000000000000",
58305 => "0000000000000000",58306 => "0000000000000000",
58307 => "0000000000000000",58308 => "0000000000000000",
58309 => "0000000000000000",58310 => "0000000000000000",
58311 => "0000000000000000",58312 => "0000000000000000",
58313 => "0000000000000000",58314 => "0000000000000000",
58315 => "0000000000000000",58316 => "0000000000000000",
58317 => "0000000000000000",58318 => "0000000000000000",
58319 => "0000000000000000",58320 => "0000000000000000",
58321 => "0000000000000000",58322 => "0000000000000000",
58323 => "0000000000000000",58324 => "0000000000000000",
58325 => "0000000000000000",58326 => "0000000000000000",
58327 => "0000000000000000",58328 => "0000000000000000",
58329 => "0000000000000000",58330 => "0000000000000000",
58331 => "0000000000000000",58332 => "0000000000000000",
58333 => "0000000000000000",58334 => "0000000000000000",
58335 => "0000000000000000",58336 => "0000000000000000",
58337 => "0000000000000000",58338 => "0000000000000000",
58339 => "0000000000000000",58340 => "0000000000000000",
58341 => "0000000000000000",58342 => "0000000000000000",
58343 => "0000000000000000",58344 => "0000000000000000",
58345 => "0000000000000000",58346 => "0000000000000000",
58347 => "0000000000000000",58348 => "0000000000000000",
58349 => "0000000000000000",58350 => "0000000000000000",
58351 => "0000000000000000",58352 => "0000000000000000",
58353 => "0000000000000000",58354 => "0000000000000000",
58355 => "0000000000000000",58356 => "0000000000000000",
58357 => "0000000000000000",58358 => "0000000000000000",
58359 => "0000000000000000",58360 => "0000000000000000",
58361 => "0000000000000000",58362 => "0000000000000000",
58363 => "0000000000000000",58364 => "0000000000000000",
58365 => "0000000000000000",58366 => "0000000000000000",
58367 => "0000000000000000",58368 => "0000000000000000",
58369 => "0000000000000000",58370 => "0000000000000000",
58371 => "0000000000000000",58372 => "0000000000000000",
58373 => "0000000000000000",58374 => "0000000000000000",
58375 => "0000000000000000",58376 => "0000000000000000",
58377 => "0000000000000000",58378 => "0000000000000000",
58379 => "0000000000000000",58380 => "0000000000000000",
58381 => "0000000000000000",58382 => "0000000000000000",
58383 => "0000000000000000",58384 => "0000000000000000",
58385 => "0000000000000000",58386 => "0000000000000000",
58387 => "0000000000000000",58388 => "0000000000000000",
58389 => "0000000000000000",58390 => "0000000000000000",
58391 => "0000000000000000",58392 => "0000000000000000",
58393 => "0000000000000000",58394 => "0000000000000000",
58395 => "0000000000000000",58396 => "0000000000000000",
58397 => "0000000000000000",58398 => "0000000000000000",
58399 => "0000000000000000",58400 => "0000000000000000",
58401 => "0000000000000000",58402 => "0000000000000000",
58403 => "0000000000000000",58404 => "0000000000000000",
58405 => "0000000000000000",58406 => "0000000000000000",
58407 => "0000000000000000",58408 => "0000000000000000",
58409 => "0000000000000000",58410 => "0000000000000000",
58411 => "0000000000000000",58412 => "0000000000000000",
58413 => "0000000000000000",58414 => "0000000000000000",
58415 => "0000000000000000",58416 => "0000000000000000",
58417 => "0000000000000000",58418 => "0000000000000000",
58419 => "0000000000000000",58420 => "0000000000000000",
58421 => "0000000000000000",58422 => "0000000000000000",
58423 => "0000000000000000",58424 => "0000000000000000",
58425 => "0000000000000000",58426 => "0000000000000000",
58427 => "0000000000000000",58428 => "0000000000000000",
58429 => "0000000000000000",58430 => "0000000000000000",
58431 => "0000000000000000",58432 => "0000000000000000",
58433 => "0000000000000000",58434 => "0000000000000000",
58435 => "0000000000000000",58436 => "0000000000000000",
58437 => "0000000000000000",58438 => "0000000000000000",
58439 => "0000000000000000",58440 => "0000000000000000",
58441 => "0000000000000000",58442 => "0000000000000000",
58443 => "0000000000000000",58444 => "0000000000000000",
58445 => "0000000000000000",58446 => "0000000000000000",
58447 => "0000000000000000",58448 => "0000000000000000",
58449 => "0000000000000000",58450 => "0000000000000000",
58451 => "0000000000000000",58452 => "0000000000000000",
58453 => "0000000000000000",58454 => "0000000000000000",
58455 => "0000000000000000",58456 => "0000000000000000",
58457 => "0000000000000000",58458 => "0000000000000000",
58459 => "0000000000000000",58460 => "0000000000000000",
58461 => "0000000000000000",58462 => "0000000000000000",
58463 => "0000000000000000",58464 => "0000000000000000",
58465 => "0000000000000000",58466 => "0000000000000000",
58467 => "0000000000000000",58468 => "0000000000000000",
58469 => "0000000000000000",58470 => "0000000000000000",
58471 => "0000000000000000",58472 => "0000000000000000",
58473 => "0000000000000000",58474 => "0000000000000000",
58475 => "0000000000000000",58476 => "0000000000000000",
58477 => "0000000000000000",58478 => "0000000000000000",
58479 => "0000000000000000",58480 => "0000000000000000",
58481 => "0000000000000000",58482 => "0000000000000000",
58483 => "0000000000000000",58484 => "0000000000000000",
58485 => "0000000000000000",58486 => "0000000000000000",
58487 => "0000000000000000",58488 => "0000000000000000",
58489 => "0000000000000000",58490 => "0000000000000000",
58491 => "0000000000000000",58492 => "0000000000000000",
58493 => "0000000000000000",58494 => "0000000000000000",
58495 => "0000000000000000",58496 => "0000000000000000",
58497 => "0000000000000000",58498 => "0000000000000000",
58499 => "0000000000000000",58500 => "0000000000000000",
58501 => "0000000000000000",58502 => "0000000000000000",
58503 => "0000000000000000",58504 => "0000000000000000",
58505 => "0000000000000000",58506 => "0000000000000000",
58507 => "0000000000000000",58508 => "0000000000000000",
58509 => "0000000000000000",58510 => "0000000000000000",
58511 => "0000000000000000",58512 => "0000000000000000",
58513 => "0000000000000000",58514 => "0000000000000000",
58515 => "0000000000000000",58516 => "0000000000000000",
58517 => "0000000000000000",58518 => "0000000000000000",
58519 => "0000000000000000",58520 => "0000000000000000",
58521 => "0000000000000000",58522 => "0000000000000000",
58523 => "0000000000000000",58524 => "0000000000000000",
58525 => "0000000000000000",58526 => "0000000000000000",
58527 => "0000000000000000",58528 => "0000000000000000",
58529 => "0000000000000000",58530 => "0000000000000000",
58531 => "0000000000000000",58532 => "0000000000000000",
58533 => "0000000000000000",58534 => "0000000000000000",
58535 => "0000000000000000",58536 => "0000000000000000",
58537 => "0000000000000000",58538 => "0000000000000000",
58539 => "0000000000000000",58540 => "0000000000000000",
58541 => "0000000000000000",58542 => "0000000000000000",
58543 => "0000000000000000",58544 => "0000000000000000",
58545 => "0000000000000000",58546 => "0000000000000000",
58547 => "0000000000000000",58548 => "0000000000000000",
58549 => "0000000000000000",58550 => "0000000000000000",
58551 => "0000000000000000",58552 => "0000000000000000",
58553 => "0000000000000000",58554 => "0000000000000000",
58555 => "0000000000000000",58556 => "0000000000000000",
58557 => "0000000000000000",58558 => "0000000000000000",
58559 => "0000000000000000",58560 => "0000000000000000",
58561 => "0000000000000000",58562 => "0000000000000000",
58563 => "0000000000000000",58564 => "0000000000000000",
58565 => "0000000000000000",58566 => "0000000000000000",
58567 => "0000000000000000",58568 => "0000000000000000",
58569 => "0000000000000000",58570 => "0000000000000000",
58571 => "0000000000000000",58572 => "0000000000000000",
58573 => "0000000000000000",58574 => "0000000000000000",
58575 => "0000000000000000",58576 => "0000000000000000",
58577 => "0000000000000000",58578 => "0000000000000000",
58579 => "0000000000000000",58580 => "0000000000000000",
58581 => "0000000000000000",58582 => "0000000000000000",
58583 => "0000000000000000",58584 => "0000000000000000",
58585 => "0000000000000000",58586 => "0000000000000000",
58587 => "0000000000000000",58588 => "0000000000000000",
58589 => "0000000000000000",58590 => "0000000000000000",
58591 => "0000000000000000",58592 => "0000000000000000",
58593 => "0000000000000000",58594 => "0000000000000000",
58595 => "0000000000000000",58596 => "0000000000000000",
58597 => "0000000000000000",58598 => "0000000000000000",
58599 => "0000000000000000",58600 => "0000000000000000",
58601 => "0000000000000000",58602 => "0000000000000000",
58603 => "0000000000000000",58604 => "0000000000000000",
58605 => "0000000000000000",58606 => "0000000000000000",
58607 => "0000000000000000",58608 => "0000000000000000",
58609 => "0000000000000000",58610 => "0000000000000000",
58611 => "0000000000000000",58612 => "0000000000000000",
58613 => "0000000000000000",58614 => "0000000000000000",
58615 => "0000000000000000",58616 => "0000000000000000",
58617 => "0000000000000000",58618 => "0000000000000000",
58619 => "0000000000000000",58620 => "0000000000000000",
58621 => "0000000000000000",58622 => "0000000000000000",
58623 => "0000000000000000",58624 => "0000000000000000",
58625 => "0000000000000000",58626 => "0000000000000000",
58627 => "0000000000000000",58628 => "0000000000000000",
58629 => "0000000000000000",58630 => "0000000000000000",
58631 => "0000000000000000",58632 => "0000000000000000",
58633 => "0000000000000000",58634 => "0000000000000000",
58635 => "0000000000000000",58636 => "0000000000000000",
58637 => "0000000000000000",58638 => "0000000000000000",
58639 => "0000000000000000",58640 => "0000000000000000",
58641 => "0000000000000000",58642 => "0000000000000000",
58643 => "0000000000000000",58644 => "0000000000000000",
58645 => "0000000000000000",58646 => "0000000000000000",
58647 => "0000000000000000",58648 => "0000000000000000",
58649 => "0000000000000000",58650 => "0000000000000000",
58651 => "0000000000000000",58652 => "0000000000000000",
58653 => "0000000000000000",58654 => "0000000000000000",
58655 => "0000000000000000",58656 => "0000000000000000",
58657 => "0000000000000000",58658 => "0000000000000000",
58659 => "0000000000000000",58660 => "0000000000000000",
58661 => "0000000000000000",58662 => "0000000000000000",
58663 => "0000000000000000",58664 => "0000000000000000",
58665 => "0000000000000000",58666 => "0000000000000000",
58667 => "0000000000000000",58668 => "0000000000000000",
58669 => "0000000000000000",58670 => "0000000000000000",
58671 => "0000000000000000",58672 => "0000000000000000",
58673 => "0000000000000000",58674 => "0000000000000000",
58675 => "0000000000000000",58676 => "0000000000000000",
58677 => "0000000000000000",58678 => "0000000000000000",
58679 => "0000000000000000",58680 => "0000000000000000",
58681 => "0000000000000000",58682 => "0000000000000000",
58683 => "0000000000000000",58684 => "0000000000000000",
58685 => "0000000000000000",58686 => "0000000000000000",
58687 => "0000000000000000",58688 => "0000000000000000",
58689 => "0000000000000000",58690 => "0000000000000000",
58691 => "0000000000000000",58692 => "0000000000000000",
58693 => "0000000000000000",58694 => "0000000000000000",
58695 => "0000000000000000",58696 => "0000000000000000",
58697 => "0000000000000000",58698 => "0000000000000000",
58699 => "0000000000000000",58700 => "0000000000000000",
58701 => "0000000000000000",58702 => "0000000000000000",
58703 => "0000000000000000",58704 => "0000000000000000",
58705 => "0000000000000000",58706 => "0000000000000000",
58707 => "0000000000000000",58708 => "0000000000000000",
58709 => "0000000000000000",58710 => "0000000000000000",
58711 => "0000000000000000",58712 => "0000000000000000",
58713 => "0000000000000000",58714 => "0000000000000000",
58715 => "0000000000000000",58716 => "0000000000000000",
58717 => "0000000000000000",58718 => "0000000000000000",
58719 => "0000000000000000",58720 => "0000000000000000",
58721 => "0000000000000000",58722 => "0000000000000000",
58723 => "0000000000000000",58724 => "0000000000000000",
58725 => "0000000000000000",58726 => "0000000000000000",
58727 => "0000000000000000",58728 => "0000000000000000",
58729 => "0000000000000000",58730 => "0000000000000000",
58731 => "0000000000000000",58732 => "0000000000000000",
58733 => "0000000000000000",58734 => "0000000000000000",
58735 => "0000000000000000",58736 => "0000000000000000",
58737 => "0000000000000000",58738 => "0000000000000000",
58739 => "0000000000000000",58740 => "0000000000000000",
58741 => "0000000000000000",58742 => "0000000000000000",
58743 => "0000000000000000",58744 => "0000000000000000",
58745 => "0000000000000000",58746 => "0000000000000000",
58747 => "0000000000000000",58748 => "0000000000000000",
58749 => "0000000000000000",58750 => "0000000000000000",
58751 => "0000000000000000",58752 => "0000000000000000",
58753 => "0000000000000000",58754 => "0000000000000000",
58755 => "0000000000000000",58756 => "0000000000000000",
58757 => "0000000000000000",58758 => "0000000000000000",
58759 => "0000000000000000",58760 => "0000000000000000",
58761 => "0000000000000000",58762 => "0000000000000000",
58763 => "0000000000000000",58764 => "0000000000000000",
58765 => "0000000000000000",58766 => "0000000000000000",
58767 => "0000000000000000",58768 => "0000000000000000",
58769 => "0000000000000000",58770 => "0000000000000000",
58771 => "0000000000000000",58772 => "0000000000000000",
58773 => "0000000000000000",58774 => "0000000000000000",
58775 => "0000000000000000",58776 => "0000000000000000",
58777 => "0000000000000000",58778 => "0000000000000000",
58779 => "0000000000000000",58780 => "0000000000000000",
58781 => "0000000000000000",58782 => "0000000000000000",
58783 => "0000000000000000",58784 => "0000000000000000",
58785 => "0000000000000000",58786 => "0000000000000000",
58787 => "0000000000000000",58788 => "0000000000000000",
58789 => "0000000000000000",58790 => "0000000000000000",
58791 => "0000000000000000",58792 => "0000000000000000",
58793 => "0000000000000000",58794 => "0000000000000000",
58795 => "0000000000000000",58796 => "0000000000000000",
58797 => "0000000000000000",58798 => "0000000000000000",
58799 => "0000000000000000",58800 => "0000000000000000",
58801 => "0000000000000000",58802 => "0000000000000000",
58803 => "0000000000000000",58804 => "0000000000000000",
58805 => "0000000000000000",58806 => "0000000000000000",
58807 => "0000000000000000",58808 => "0000000000000000",
58809 => "0000000000000000",58810 => "0000000000000000",
58811 => "0000000000000000",58812 => "0000000000000000",
58813 => "0000000000000000",58814 => "0000000000000000",
58815 => "0000000000000000",58816 => "0000000000000000",
58817 => "0000000000000000",58818 => "0000000000000000",
58819 => "0000000000000000",58820 => "0000000000000000",
58821 => "0000000000000000",58822 => "0000000000000000",
58823 => "0000000000000000",58824 => "0000000000000000",
58825 => "0000000000000000",58826 => "0000000000000000",
58827 => "0000000000000000",58828 => "0000000000000000",
58829 => "0000000000000000",58830 => "0000000000000000",
58831 => "0000000000000000",58832 => "0000000000000000",
58833 => "0000000000000000",58834 => "0000000000000000",
58835 => "0000000000000000",58836 => "0000000000000000",
58837 => "0000000000000000",58838 => "0000000000000000",
58839 => "0000000000000000",58840 => "0000000000000000",
58841 => "0000000000000000",58842 => "0000000000000000",
58843 => "0000000000000000",58844 => "0000000000000000",
58845 => "0000000000000000",58846 => "0000000000000000",
58847 => "0000000000000000",58848 => "0000000000000000",
58849 => "0000000000000000",58850 => "0000000000000000",
58851 => "0000000000000000",58852 => "0000000000000000",
58853 => "0000000000000000",58854 => "0000000000000000",
58855 => "0000000000000000",58856 => "0000000000000000",
58857 => "0000000000000000",58858 => "0000000000000000",
58859 => "0000000000000000",58860 => "0000000000000000",
58861 => "0000000000000000",58862 => "0000000000000000",
58863 => "0000000000000000",58864 => "0000000000000000",
58865 => "0000000000000000",58866 => "0000000000000000",
58867 => "0000000000000000",58868 => "0000000000000000",
58869 => "0000000000000000",58870 => "0000000000000000",
58871 => "0000000000000000",58872 => "0000000000000000",
58873 => "0000000000000000",58874 => "0000000000000000",
58875 => "0000000000000000",58876 => "0000000000000000",
58877 => "0000000000000000",58878 => "0000000000000000",
58879 => "0000000000000000",58880 => "0000000000000000",
58881 => "0000000000000000",58882 => "0000000000000000",
58883 => "0000000000000000",58884 => "0000000000000000",
58885 => "0000000000000000",58886 => "0000000000000000",
58887 => "0000000000000000",58888 => "0000000000000000",
58889 => "0000000000000000",58890 => "0000000000000000",
58891 => "0000000000000000",58892 => "0000000000000000",
58893 => "0000000000000000",58894 => "0000000000000000",
58895 => "0000000000000000",58896 => "0000000000000000",
58897 => "0000000000000000",58898 => "0000000000000000",
58899 => "0000000000000000",58900 => "0000000000000000",
58901 => "0000000000000000",58902 => "0000000000000000",
58903 => "0000000000000000",58904 => "0000000000000000",
58905 => "0000000000000000",58906 => "0000000000000000",
58907 => "0000000000000000",58908 => "0000000000000000",
58909 => "0000000000000000",58910 => "0000000000000000",
58911 => "0000000000000000",58912 => "0000000000000000",
58913 => "0000000000000000",58914 => "0000000000000000",
58915 => "0000000000000000",58916 => "0000000000000000",
58917 => "0000000000000000",58918 => "0000000000000000",
58919 => "0000000000000000",58920 => "0000000000000000",
58921 => "0000000000000000",58922 => "0000000000000000",
58923 => "0000000000000000",58924 => "0000000000000000",
58925 => "0000000000000000",58926 => "0000000000000000",
58927 => "0000000000000000",58928 => "0000000000000000",
58929 => "0000000000000000",58930 => "0000000000000000",
58931 => "0000000000000000",58932 => "0000000000000000",
58933 => "0000000000000000",58934 => "0000000000000000",
58935 => "0000000000000000",58936 => "0000000000000000",
58937 => "0000000000000000",58938 => "0000000000000000",
58939 => "0000000000000000",58940 => "0000000000000000",
58941 => "0000000000000000",58942 => "0000000000000000",
58943 => "0000000000000000",58944 => "0000000000000000",
58945 => "0000000000000000",58946 => "0000000000000000",
58947 => "0000000000000000",58948 => "0000000000000000",
58949 => "0000000000000000",58950 => "0000000000000000",
58951 => "0000000000000000",58952 => "0000000000000000",
58953 => "0000000000000000",58954 => "0000000000000000",
58955 => "0000000000000000",58956 => "0000000000000000",
58957 => "0000000000000000",58958 => "0000000000000000",
58959 => "0000000000000000",58960 => "0000000000000000",
58961 => "0000000000000000",58962 => "0000000000000000",
58963 => "0000000000000000",58964 => "0000000000000000",
58965 => "0000000000000000",58966 => "0000000000000000",
58967 => "0000000000000000",58968 => "0000000000000000",
58969 => "0000000000000000",58970 => "0000000000000000",
58971 => "0000000000000000",58972 => "0000000000000000",
58973 => "0000000000000000",58974 => "0000000000000000",
58975 => "0000000000000000",58976 => "0000000000000000",
58977 => "0000000000000000",58978 => "0000000000000000",
58979 => "0000000000000000",58980 => "0000000000000000",
58981 => "0000000000000000",58982 => "0000000000000000",
58983 => "0000000000000000",58984 => "0000000000000000",
58985 => "0000000000000000",58986 => "0000000000000000",
58987 => "0000000000000000",58988 => "0000000000000000",
58989 => "0000000000000000",58990 => "0000000000000000",
58991 => "0000000000000000",58992 => "0000000000000000",
58993 => "0000000000000000",58994 => "0000000000000000",
58995 => "0000000000000000",58996 => "0000000000000000",
58997 => "0000000000000000",58998 => "0000000000000000",
58999 => "0000000000000000",59000 => "0000000000000000",
59001 => "0000000000000000",59002 => "0000000000000000",
59003 => "0000000000000000",59004 => "0000000000000000",
59005 => "0000000000000000",59006 => "0000000000000000",
59007 => "0000000000000000",59008 => "0000000000000000",
59009 => "0000000000000000",59010 => "0000000000000000",
59011 => "0000000000000000",59012 => "0000000000000000",
59013 => "0000000000000000",59014 => "0000000000000000",
59015 => "0000000000000000",59016 => "0000000000000000",
59017 => "0000000000000000",59018 => "0000000000000000",
59019 => "0000000000000000",59020 => "0000000000000000",
59021 => "0000000000000000",59022 => "0000000000000000",
59023 => "0000000000000000",59024 => "0000000000000000",
59025 => "0000000000000000",59026 => "0000000000000000",
59027 => "0000000000000000",59028 => "0000000000000000",
59029 => "0000000000000000",59030 => "0000000000000000",
59031 => "0000000000000000",59032 => "0000000000000000",
59033 => "0000000000000000",59034 => "0000000000000000",
59035 => "0000000000000000",59036 => "0000000000000000",
59037 => "0000000000000000",59038 => "0000000000000000",
59039 => "0000000000000000",59040 => "0000000000000000",
59041 => "0000000000000000",59042 => "0000000000000000",
59043 => "0000000000000000",59044 => "0000000000000000",
59045 => "0000000000000000",59046 => "0000000000000000",
59047 => "0000000000000000",59048 => "0000000000000000",
59049 => "0000000000000000",59050 => "0000000000000000",
59051 => "0000000000000000",59052 => "0000000000000000",
59053 => "0000000000000000",59054 => "0000000000000000",
59055 => "0000000000000000",59056 => "0000000000000000",
59057 => "0000000000000000",59058 => "0000000000000000",
59059 => "0000000000000000",59060 => "0000000000000000",
59061 => "0000000000000000",59062 => "0000000000000000",
59063 => "0000000000000000",59064 => "0000000000000000",
59065 => "0000000000000000",59066 => "0000000000000000",
59067 => "0000000000000000",59068 => "0000000000000000",
59069 => "0000000000000000",59070 => "0000000000000000",
59071 => "0000000000000000",59072 => "0000000000000000",
59073 => "0000000000000000",59074 => "0000000000000000",
59075 => "0000000000000000",59076 => "0000000000000000",
59077 => "0000000000000000",59078 => "0000000000000000",
59079 => "0000000000000000",59080 => "0000000000000000",
59081 => "0000000000000000",59082 => "0000000000000000",
59083 => "0000000000000000",59084 => "0000000000000000",
59085 => "0000000000000000",59086 => "0000000000000000",
59087 => "0000000000000000",59088 => "0000000000000000",
59089 => "0000000000000000",59090 => "0000000000000000",
59091 => "0000000000000000",59092 => "0000000000000000",
59093 => "0000000000000000",59094 => "0000000000000000",
59095 => "0000000000000000",59096 => "0000000000000000",
59097 => "0000000000000000",59098 => "0000000000000000",
59099 => "0000000000000000",59100 => "0000000000000000",
59101 => "0000000000000000",59102 => "0000000000000000",
59103 => "0000000000000000",59104 => "0000000000000000",
59105 => "0000000000000000",59106 => "0000000000000000",
59107 => "0000000000000000",59108 => "0000000000000000",
59109 => "0000000000000000",59110 => "0000000000000000",
59111 => "0000000000000000",59112 => "0000000000000000",
59113 => "0000000000000000",59114 => "0000000000000000",
59115 => "0000000000000000",59116 => "0000000000000000",
59117 => "0000000000000000",59118 => "0000000000000000",
59119 => "0000000000000000",59120 => "0000000000000000",
59121 => "0000000000000000",59122 => "0000000000000000",
59123 => "0000000000000000",59124 => "0000000000000000",
59125 => "0000000000000000",59126 => "0000000000000000",
59127 => "0000000000000000",59128 => "0000000000000000",
59129 => "0000000000000000",59130 => "0000000000000000",
59131 => "0000000000000000",59132 => "0000000000000000",
59133 => "0000000000000000",59134 => "0000000000000000",
59135 => "0000000000000000",59136 => "0000000000000000",
59137 => "0000000000000000",59138 => "0000000000000000",
59139 => "0000000000000000",59140 => "0000000000000000",
59141 => "0000000000000000",59142 => "0000000000000000",
59143 => "0000000000000000",59144 => "0000000000000000",
59145 => "0000000000000000",59146 => "0000000000000000",
59147 => "0000000000000000",59148 => "0000000000000000",
59149 => "0000000000000000",59150 => "0000000000000000",
59151 => "0000000000000000",59152 => "0000000000000000",
59153 => "0000000000000000",59154 => "0000000000000000",
59155 => "0000000000000000",59156 => "0000000000000000",
59157 => "0000000000000000",59158 => "0000000000000000",
59159 => "0000000000000000",59160 => "0000000000000000",
59161 => "0000000000000000",59162 => "0000000000000000",
59163 => "0000000000000000",59164 => "0000000000000000",
59165 => "0000000000000000",59166 => "0000000000000000",
59167 => "0000000000000000",59168 => "0000000000000000",
59169 => "0000000000000000",59170 => "0000000000000000",
59171 => "0000000000000000",59172 => "0000000000000000",
59173 => "0000000000000000",59174 => "0000000000000000",
59175 => "0000000000000000",59176 => "0000000000000000",
59177 => "0000000000000000",59178 => "0000000000000000",
59179 => "0000000000000000",59180 => "0000000000000000",
59181 => "0000000000000000",59182 => "0000000000000000",
59183 => "0000000000000000",59184 => "0000000000000000",
59185 => "0000000000000000",59186 => "0000000000000000",
59187 => "0000000000000000",59188 => "0000000000000000",
59189 => "0000000000000000",59190 => "0000000000000000",
59191 => "0000000000000000",59192 => "0000000000000000",
59193 => "0000000000000000",59194 => "0000000000000000",
59195 => "0000000000000000",59196 => "0000000000000000",
59197 => "0000000000000000",59198 => "0000000000000000",
59199 => "0000000000000000",59200 => "0000000000000000",
59201 => "0000000000000000",59202 => "0000000000000000",
59203 => "0000000000000000",59204 => "0000000000000000",
59205 => "0000000000000000",59206 => "0000000000000000",
59207 => "0000000000000000",59208 => "0000000000000000",
59209 => "0000000000000000",59210 => "0000000000000000",
59211 => "0000000000000000",59212 => "0000000000000000",
59213 => "0000000000000000",59214 => "0000000000000000",
59215 => "0000000000000000",59216 => "0000000000000000",
59217 => "0000000000000000",59218 => "0000000000000000",
59219 => "0000000000000000",59220 => "0000000000000000",
59221 => "0000000000000000",59222 => "0000000000000000",
59223 => "0000000000000000",59224 => "0000000000000000",
59225 => "0000000000000000",59226 => "0000000000000000",
59227 => "0000000000000000",59228 => "0000000000000000",
59229 => "0000000000000000",59230 => "0000000000000000",
59231 => "0000000000000000",59232 => "0000000000000000",
59233 => "0000000000000000",59234 => "0000000000000000",
59235 => "0000000000000000",59236 => "0000000000000000",
59237 => "0000000000000000",59238 => "0000000000000000",
59239 => "0000000000000000",59240 => "0000000000000000",
59241 => "0000000000000000",59242 => "0000000000000000",
59243 => "0000000000000000",59244 => "0000000000000000",
59245 => "0000000000000000",59246 => "0000000000000000",
59247 => "0000000000000000",59248 => "0000000000000000",
59249 => "0000000000000000",59250 => "0000000000000000",
59251 => "0000000000000000",59252 => "0000000000000000",
59253 => "0000000000000000",59254 => "0000000000000000",
59255 => "0000000000000000",59256 => "0000000000000000",
59257 => "0000000000000000",59258 => "0000000000000000",
59259 => "0000000000000000",59260 => "0000000000000000",
59261 => "0000000000000000",59262 => "0000000000000000",
59263 => "0000000000000000",59264 => "0000000000000000",
59265 => "0000000000000000",59266 => "0000000000000000",
59267 => "0000000000000000",59268 => "0000000000000000",
59269 => "0000000000000000",59270 => "0000000000000000",
59271 => "0000000000000000",59272 => "0000000000000000",
59273 => "0000000000000000",59274 => "0000000000000000",
59275 => "0000000000000000",59276 => "0000000000000000",
59277 => "0000000000000000",59278 => "0000000000000000",
59279 => "0000000000000000",59280 => "0000000000000000",
59281 => "0000000000000000",59282 => "0000000000000000",
59283 => "0000000000000000",59284 => "0000000000000000",
59285 => "0000000000000000",59286 => "0000000000000000",
59287 => "0000000000000000",59288 => "0000000000000000",
59289 => "0000000000000000",59290 => "0000000000000000",
59291 => "0000000000000000",59292 => "0000000000000000",
59293 => "0000000000000000",59294 => "0000000000000000",
59295 => "0000000000000000",59296 => "0000000000000000",
59297 => "0000000000000000",59298 => "0000000000000000",
59299 => "0000000000000000",59300 => "0000000000000000",
59301 => "0000000000000000",59302 => "0000000000000000",
59303 => "0000000000000000",59304 => "0000000000000000",
59305 => "0000000000000000",59306 => "0000000000000000",
59307 => "0000000000000000",59308 => "0000000000000000",
59309 => "0000000000000000",59310 => "0000000000000000",
59311 => "0000000000000000",59312 => "0000000000000000",
59313 => "0000000000000000",59314 => "0000000000000000",
59315 => "0000000000000000",59316 => "0000000000000000",
59317 => "0000000000000000",59318 => "0000000000000000",
59319 => "0000000000000000",59320 => "0000000000000000",
59321 => "0000000000000000",59322 => "0000000000000000",
59323 => "0000000000000000",59324 => "0000000000000000",
59325 => "0000000000000000",59326 => "0000000000000000",
59327 => "0000000000000000",59328 => "0000000000000000",
59329 => "0000000000000000",59330 => "0000000000000000",
59331 => "0000000000000000",59332 => "0000000000000000",
59333 => "0000000000000000",59334 => "0000000000000000",
59335 => "0000000000000000",59336 => "0000000000000000",
59337 => "0000000000000000",59338 => "0000000000000000",
59339 => "0000000000000000",59340 => "0000000000000000",
59341 => "0000000000000000",59342 => "0000000000000000",
59343 => "0000000000000000",59344 => "0000000000000000",
59345 => "0000000000000000",59346 => "0000000000000000",
59347 => "0000000000000000",59348 => "0000000000000000",
59349 => "0000000000000000",59350 => "0000000000000000",
59351 => "0000000000000000",59352 => "0000000000000000",
59353 => "0000000000000000",59354 => "0000000000000000",
59355 => "0000000000000000",59356 => "0000000000000000",
59357 => "0000000000000000",59358 => "0000000000000000",
59359 => "0000000000000000",59360 => "0000000000000000",
59361 => "0000000000000000",59362 => "0000000000000000",
59363 => "0000000000000000",59364 => "0000000000000000",
59365 => "0000000000000000",59366 => "0000000000000000",
59367 => "0000000000000000",59368 => "0000000000000000",
59369 => "0000000000000000",59370 => "0000000000000000",
59371 => "0000000000000000",59372 => "0000000000000000",
59373 => "0000000000000000",59374 => "0000000000000000",
59375 => "0000000000000000",59376 => "0000000000000000",
59377 => "0000000000000000",59378 => "0000000000000000",
59379 => "0000000000000000",59380 => "0000000000000000",
59381 => "0000000000000000",59382 => "0000000000000000",
59383 => "0000000000000000",59384 => "0000000000000000",
59385 => "0000000000000000",59386 => "0000000000000000",
59387 => "0000000000000000",59388 => "0000000000000000",
59389 => "0000000000000000",59390 => "0000000000000000",
59391 => "0000000000000000",59392 => "0000000000000000",
59393 => "0000000000000000",59394 => "0000000000000000",
59395 => "0000000000000000",59396 => "0000000000000000",
59397 => "0000000000000000",59398 => "0000000000000000",
59399 => "0000000000000000",59400 => "0000000000000000",
59401 => "0000000000000000",59402 => "0000000000000000",
59403 => "0000000000000000",59404 => "0000000000000000",
59405 => "0000000000000000",59406 => "0000000000000000",
59407 => "0000000000000000",59408 => "0000000000000000",
59409 => "0000000000000000",59410 => "0000000000000000",
59411 => "0000000000000000",59412 => "0000000000000000",
59413 => "0000000000000000",59414 => "0000000000000000",
59415 => "0000000000000000",59416 => "0000000000000000",
59417 => "0000000000000000",59418 => "0000000000000000",
59419 => "0000000000000000",59420 => "0000000000000000",
59421 => "0000000000000000",59422 => "0000000000000000",
59423 => "0000000000000000",59424 => "0000000000000000",
59425 => "0000000000000000",59426 => "0000000000000000",
59427 => "0000000000000000",59428 => "0000000000000000",
59429 => "0000000000000000",59430 => "0000000000000000",
59431 => "0000000000000000",59432 => "0000000000000000",
59433 => "0000000000000000",59434 => "0000000000000000",
59435 => "0000000000000000",59436 => "0000000000000000",
59437 => "0000000000000000",59438 => "0000000000000000",
59439 => "0000000000000000",59440 => "0000000000000000",
59441 => "0000000000000000",59442 => "0000000000000000",
59443 => "0000000000000000",59444 => "0000000000000000",
59445 => "0000000000000000",59446 => "0000000000000000",
59447 => "0000000000000000",59448 => "0000000000000000",
59449 => "0000000000000000",59450 => "0000000000000000",
59451 => "0000000000000000",59452 => "0000000000000000",
59453 => "0000000000000000",59454 => "0000000000000000",
59455 => "0000000000000000",59456 => "0000000000000000",
59457 => "0000000000000000",59458 => "0000000000000000",
59459 => "0000000000000000",59460 => "0000000000000000",
59461 => "0000000000000000",59462 => "0000000000000000",
59463 => "0000000000000000",59464 => "0000000000000000",
59465 => "0000000000000000",59466 => "0000000000000000",
59467 => "0000000000000000",59468 => "0000000000000000",
59469 => "0000000000000000",59470 => "0000000000000000",
59471 => "0000000000000000",59472 => "0000000000000000",
59473 => "0000000000000000",59474 => "0000000000000000",
59475 => "0000000000000000",59476 => "0000000000000000",
59477 => "0000000000000000",59478 => "0000000000000000",
59479 => "0000000000000000",59480 => "0000000000000000",
59481 => "0000000000000000",59482 => "0000000000000000",
59483 => "0000000000000000",59484 => "0000000000000000",
59485 => "0000000000000000",59486 => "0000000000000000",
59487 => "0000000000000000",59488 => "0000000000000000",
59489 => "0000000000000000",59490 => "0000000000000000",
59491 => "0000000000000000",59492 => "0000000000000000",
59493 => "0000000000000000",59494 => "0000000000000000",
59495 => "0000000000000000",59496 => "0000000000000000",
59497 => "0000000000000000",59498 => "0000000000000000",
59499 => "0000000000000000",59500 => "0000000000000000",
59501 => "0000000000000000",59502 => "0000000000000000",
59503 => "0000000000000000",59504 => "0000000000000000",
59505 => "0000000000000000",59506 => "0000000000000000",
59507 => "0000000000000000",59508 => "0000000000000000",
59509 => "0000000000000000",59510 => "0000000000000000",
59511 => "0000000000000000",59512 => "0000000000000000",
59513 => "0000000000000000",59514 => "0000000000000000",
59515 => "0000000000000000",59516 => "0000000000000000",
59517 => "0000000000000000",59518 => "0000000000000000",
59519 => "0000000000000000",59520 => "0000000000000000",
59521 => "0000000000000000",59522 => "0000000000000000",
59523 => "0000000000000000",59524 => "0000000000000000",
59525 => "0000000000000000",59526 => "0000000000000000",
59527 => "0000000000000000",59528 => "0000000000000000",
59529 => "0000000000000000",59530 => "0000000000000000",
59531 => "0000000000000000",59532 => "0000000000000000",
59533 => "0000000000000000",59534 => "0000000000000000",
59535 => "0000000000000000",59536 => "0000000000000000",
59537 => "0000000000000000",59538 => "0000000000000000",
59539 => "0000000000000000",59540 => "0000000000000000",
59541 => "0000000000000000",59542 => "0000000000000000",
59543 => "0000000000000000",59544 => "0000000000000000",
59545 => "0000000000000000",59546 => "0000000000000000",
59547 => "0000000000000000",59548 => "0000000000000000",
59549 => "0000000000000000",59550 => "0000000000000000",
59551 => "0000000000000000",59552 => "0000000000000000",
59553 => "0000000000000000",59554 => "0000000000000000",
59555 => "0000000000000000",59556 => "0000000000000000",
59557 => "0000000000000000",59558 => "0000000000000000",
59559 => "0000000000000000",59560 => "0000000000000000",
59561 => "0000000000000000",59562 => "0000000000000000",
59563 => "0000000000000000",59564 => "0000000000000000",
59565 => "0000000000000000",59566 => "0000000000000000",
59567 => "0000000000000000",59568 => "0000000000000000",
59569 => "0000000000000000",59570 => "0000000000000000",
59571 => "0000000000000000",59572 => "0000000000000000",
59573 => "0000000000000000",59574 => "0000000000000000",
59575 => "0000000000000000",59576 => "0000000000000000",
59577 => "0000000000000000",59578 => "0000000000000000",
59579 => "0000000000000000",59580 => "0000000000000000",
59581 => "0000000000000000",59582 => "0000000000000000",
59583 => "0000000000000000",59584 => "0000000000000000",
59585 => "0000000000000000",59586 => "0000000000000000",
59587 => "0000000000000000",59588 => "0000000000000000",
59589 => "0000000000000000",59590 => "0000000000000000",
59591 => "0000000000000000",59592 => "0000000000000000",
59593 => "0000000000000000",59594 => "0000000000000000",
59595 => "0000000000000000",59596 => "0000000000000000",
59597 => "0000000000000000",59598 => "0000000000000000",
59599 => "0000000000000000",59600 => "0000000000000000",
59601 => "0000000000000000",59602 => "0000000000000000",
59603 => "0000000000000000",59604 => "0000000000000000",
59605 => "0000000000000000",59606 => "0000000000000000",
59607 => "0000000000000000",59608 => "0000000000000000",
59609 => "0000000000000000",59610 => "0000000000000000",
59611 => "0000000000000000",59612 => "0000000000000000",
59613 => "0000000000000000",59614 => "0000000000000000",
59615 => "0000000000000000",59616 => "0000000000000000",
59617 => "0000000000000000",59618 => "0000000000000000",
59619 => "0000000000000000",59620 => "0000000000000000",
59621 => "0000000000000000",59622 => "0000000000000000",
59623 => "0000000000000000",59624 => "0000000000000000",
59625 => "0000000000000000",59626 => "0000000000000000",
59627 => "0000000000000000",59628 => "0000000000000000",
59629 => "0000000000000000",59630 => "0000000000000000",
59631 => "0000000000000000",59632 => "0000000000000000",
59633 => "0000000000000000",59634 => "0000000000000000",
59635 => "0000000000000000",59636 => "0000000000000000",
59637 => "0000000000000000",59638 => "0000000000000000",
59639 => "0000000000000000",59640 => "0000000000000000",
59641 => "0000000000000000",59642 => "0000000000000000",
59643 => "0000000000000000",59644 => "0000000000000000",
59645 => "0000000000000000",59646 => "0000000000000000",
59647 => "0000000000000000",59648 => "0000000000000000",
59649 => "0000000000000000",59650 => "0000000000000000",
59651 => "0000000000000000",59652 => "0000000000000000",
59653 => "0000000000000000",59654 => "0000000000000000",
59655 => "0000000000000000",59656 => "0000000000000000",
59657 => "0000000000000000",59658 => "0000000000000000",
59659 => "0000000000000000",59660 => "0000000000000000",
59661 => "0000000000000000",59662 => "0000000000000000",
59663 => "0000000000000000",59664 => "0000000000000000",
59665 => "0000000000000000",59666 => "0000000000000000",
59667 => "0000000000000000",59668 => "0000000000000000",
59669 => "0000000000000000",59670 => "0000000000000000",
59671 => "0000000000000000",59672 => "0000000000000000",
59673 => "0000000000000000",59674 => "0000000000000000",
59675 => "0000000000000000",59676 => "0000000000000000",
59677 => "0000000000000000",59678 => "0000000000000000",
59679 => "0000000000000000",59680 => "0000000000000000",
59681 => "0000000000000000",59682 => "0000000000000000",
59683 => "0000000000000000",59684 => "0000000000000000",
59685 => "0000000000000000",59686 => "0000000000000000",
59687 => "0000000000000000",59688 => "0000000000000000",
59689 => "0000000000000000",59690 => "0000000000000000",
59691 => "0000000000000000",59692 => "0000000000000000",
59693 => "0000000000000000",59694 => "0000000000000000",
59695 => "0000000000000000",59696 => "0000000000000000",
59697 => "0000000000000000",59698 => "0000000000000000",
59699 => "0000000000000000",59700 => "0000000000000000",
59701 => "0000000000000000",59702 => "0000000000000000",
59703 => "0000000000000000",59704 => "0000000000000000",
59705 => "0000000000000000",59706 => "0000000000000000",
59707 => "0000000000000000",59708 => "0000000000000000",
59709 => "0000000000000000",59710 => "0000000000000000",
59711 => "0000000000000000",59712 => "0000000000000000",
59713 => "0000000000000000",59714 => "0000000000000000",
59715 => "0000000000000000",59716 => "0000000000000000",
59717 => "0000000000000000",59718 => "0000000000000000",
59719 => "0000000000000000",59720 => "0000000000000000",
59721 => "0000000000000000",59722 => "0000000000000000",
59723 => "0000000000000000",59724 => "0000000000000000",
59725 => "0000000000000000",59726 => "0000000000000000",
59727 => "0000000000000000",59728 => "0000000000000000",
59729 => "0000000000000000",59730 => "0000000000000000",
59731 => "0000000000000000",59732 => "0000000000000000",
59733 => "0000000000000000",59734 => "0000000000000000",
59735 => "0000000000000000",59736 => "0000000000000000",
59737 => "0000000000000000",59738 => "0000000000000000",
59739 => "0000000000000000",59740 => "0000000000000000",
59741 => "0000000000000000",59742 => "0000000000000000",
59743 => "0000000000000000",59744 => "0000000000000000",
59745 => "0000000000000000",59746 => "0000000000000000",
59747 => "0000000000000000",59748 => "0000000000000000",
59749 => "0000000000000000",59750 => "0000000000000000",
59751 => "0000000000000000",59752 => "0000000000000000",
59753 => "0000000000000000",59754 => "0000000000000000",
59755 => "0000000000000000",59756 => "0000000000000000",
59757 => "0000000000000000",59758 => "0000000000000000",
59759 => "0000000000000000",59760 => "0000000000000000",
59761 => "0000000000000000",59762 => "0000000000000000",
59763 => "0000000000000000",59764 => "0000000000000000",
59765 => "0000000000000000",59766 => "0000000000000000",
59767 => "0000000000000000",59768 => "0000000000000000",
59769 => "0000000000000000",59770 => "0000000000000000",
59771 => "0000000000000000",59772 => "0000000000000000",
59773 => "0000000000000000",59774 => "0000000000000000",
59775 => "0000000000000000",59776 => "0000000000000000",
59777 => "0000000000000000",59778 => "0000000000000000",
59779 => "0000000000000000",59780 => "0000000000000000",
59781 => "0000000000000000",59782 => "0000000000000000",
59783 => "0000000000000000",59784 => "0000000000000000",
59785 => "0000000000000000",59786 => "0000000000000000",
59787 => "0000000000000000",59788 => "0000000000000000",
59789 => "0000000000000000",59790 => "0000000000000000",
59791 => "0000000000000000",59792 => "0000000000000000",
59793 => "0000000000000000",59794 => "0000000000000000",
59795 => "0000000000000000",59796 => "0000000000000000",
59797 => "0000000000000000",59798 => "0000000000000000",
59799 => "0000000000000000",59800 => "0000000000000000",
59801 => "0000000000000000",59802 => "0000000000000000",
59803 => "0000000000000000",59804 => "0000000000000000",
59805 => "0000000000000000",59806 => "0000000000000000",
59807 => "0000000000000000",59808 => "0000000000000000",
59809 => "0000000000000000",59810 => "0000000000000000",
59811 => "0000000000000000",59812 => "0000000000000000",
59813 => "0000000000000000",59814 => "0000000000000000",
59815 => "0000000000000000",59816 => "0000000000000000",
59817 => "0000000000000000",59818 => "0000000000000000",
59819 => "0000000000000000",59820 => "0000000000000000",
59821 => "0000000000000000",59822 => "0000000000000000",
59823 => "0000000000000000",59824 => "0000000000000000",
59825 => "0000000000000000",59826 => "0000000000000000",
59827 => "0000000000000000",59828 => "0000000000000000",
59829 => "0000000000000000",59830 => "0000000000000000",
59831 => "0000000000000000",59832 => "0000000000000000",
59833 => "0000000000000000",59834 => "0000000000000000",
59835 => "0000000000000000",59836 => "0000000000000000",
59837 => "0000000000000000",59838 => "0000000000000000",
59839 => "0000000000000000",59840 => "0000000000000000",
59841 => "0000000000000000",59842 => "0000000000000000",
59843 => "0000000000000000",59844 => "0000000000000000",
59845 => "0000000000000000",59846 => "0000000000000000",
59847 => "0000000000000000",59848 => "0000000000000000",
59849 => "0000000000000000",59850 => "0000000000000000",
59851 => "0000000000000000",59852 => "0000000000000000",
59853 => "0000000000000000",59854 => "0000000000000000",
59855 => "0000000000000000",59856 => "0000000000000000",
59857 => "0000000000000000",59858 => "0000000000000000",
59859 => "0000000000000000",59860 => "0000000000000000",
59861 => "0000000000000000",59862 => "0000000000000000",
59863 => "0000000000000000",59864 => "0000000000000000",
59865 => "0000000000000000",59866 => "0000000000000000",
59867 => "0000000000000000",59868 => "0000000000000000",
59869 => "0000000000000000",59870 => "0000000000000000",
59871 => "0000000000000000",59872 => "0000000000000000",
59873 => "0000000000000000",59874 => "0000000000000000",
59875 => "0000000000000000",59876 => "0000000000000000",
59877 => "0000000000000000",59878 => "0000000000000000",
59879 => "0000000000000000",59880 => "0000000000000000",
59881 => "0000000000000000",59882 => "0000000000000000",
59883 => "0000000000000000",59884 => "0000000000000000",
59885 => "0000000000000000",59886 => "0000000000000000",
59887 => "0000000000000000",59888 => "0000000000000000",
59889 => "0000000000000000",59890 => "0000000000000000",
59891 => "0000000000000000",59892 => "0000000000000000",
59893 => "0000000000000000",59894 => "0000000000000000",
59895 => "0000000000000000",59896 => "0000000000000000",
59897 => "0000000000000000",59898 => "0000000000000000",
59899 => "0000000000000000",59900 => "0000000000000000",
59901 => "0000000000000000",59902 => "0000000000000000",
59903 => "0000000000000000",59904 => "0000000000000000",
59905 => "0000000000000000",59906 => "0000000000000000",
59907 => "0000000000000000",59908 => "0000000000000000",
59909 => "0000000000000000",59910 => "0000000000000000",
59911 => "0000000000000000",59912 => "0000000000000000",
59913 => "0000000000000000",59914 => "0000000000000000",
59915 => "0000000000000000",59916 => "0000000000000000",
59917 => "0000000000000000",59918 => "0000000000000000",
59919 => "0000000000000000",59920 => "0000000000000000",
59921 => "0000000000000000",59922 => "0000000000000000",
59923 => "0000000000000000",59924 => "0000000000000000",
59925 => "0000000000000000",59926 => "0000000000000000",
59927 => "0000000000000000",59928 => "0000000000000000",
59929 => "0000000000000000",59930 => "0000000000000000",
59931 => "0000000000000000",59932 => "0000000000000000",
59933 => "0000000000000000",59934 => "0000000000000000",
59935 => "0000000000000000",59936 => "0000000000000000",
59937 => "0000000000000000",59938 => "0000000000000000",
59939 => "0000000000000000",59940 => "0000000000000000",
59941 => "0000000000000000",59942 => "0000000000000000",
59943 => "0000000000000000",59944 => "0000000000000000",
59945 => "0000000000000000",59946 => "0000000000000000",
59947 => "0000000000000000",59948 => "0000000000000000",
59949 => "0000000000000000",59950 => "0000000000000000",
59951 => "0000000000000000",59952 => "0000000000000000",
59953 => "0000000000000000",59954 => "0000000000000000",
59955 => "0000000000000000",59956 => "0000000000000000",
59957 => "0000000000000000",59958 => "0000000000000000",
59959 => "0000000000000000",59960 => "0000000000000000",
59961 => "0000000000000000",59962 => "0000000000000000",
59963 => "0000000000000000",59964 => "0000000000000000",
59965 => "0000000000000000",59966 => "0000000000000000",
59967 => "0000000000000000",59968 => "0000000000000000",
59969 => "0000000000000000",59970 => "0000000000000000",
59971 => "0000000000000000",59972 => "0000000000000000",
59973 => "0000000000000000",59974 => "0000000000000000",
59975 => "0000000000000000",59976 => "0000000000000000",
59977 => "0000000000000000",59978 => "0000000000000000",
59979 => "0000000000000000",59980 => "0000000000000000",
59981 => "0000000000000000",59982 => "0000000000000000",
59983 => "0000000000000000",59984 => "0000000000000000",
59985 => "0000000000000000",59986 => "0000000000000000",
59987 => "0000000000000000",59988 => "0000000000000000",
59989 => "0000000000000000",59990 => "0000000000000000",
59991 => "0000000000000000",59992 => "0000000000000000",
59993 => "0000000000000000",59994 => "0000000000000000",
59995 => "0000000000000000",59996 => "0000000000000000",
59997 => "0000000000000000",59998 => "0000000000000000",
59999 => "0000000000000000",60000 => "0000000000000000",
60001 => "0000000000000000",60002 => "0000000000000000",
60003 => "0000000000000000",60004 => "0000000000000000",
60005 => "0000000000000000",60006 => "0000000000000000",
60007 => "0000000000000000",60008 => "0000000000000000",
60009 => "0000000000000000",60010 => "0000000000000000",
60011 => "0000000000000000",60012 => "0000000000000000",
60013 => "0000000000000000",60014 => "0000000000000000",
60015 => "0000000000000000",60016 => "0000000000000000",
60017 => "0000000000000000",60018 => "0000000000000000",
60019 => "0000000000000000",60020 => "0000000000000000",
60021 => "0000000000000000",60022 => "0000000000000000",
60023 => "0000000000000000",60024 => "0000000000000000",
60025 => "0000000000000000",60026 => "0000000000000000",
60027 => "0000000000000000",60028 => "0000000000000000",
60029 => "0000000000000000",60030 => "0000000000000000",
60031 => "0000000000000000",60032 => "0000000000000000",
60033 => "0000000000000000",60034 => "0000000000000000",
60035 => "0000000000000000",60036 => "0000000000000000",
60037 => "0000000000000000",60038 => "0000000000000000",
60039 => "0000000000000000",60040 => "0000000000000000",
60041 => "0000000000000000",60042 => "0000000000000000",
60043 => "0000000000000000",60044 => "0000000000000000",
60045 => "0000000000000000",60046 => "0000000000000000",
60047 => "0000000000000000",60048 => "0000000000000000",
60049 => "0000000000000000",60050 => "0000000000000000",
60051 => "0000000000000000",60052 => "0000000000000000",
60053 => "0000000000000000",60054 => "0000000000000000",
60055 => "0000000000000000",60056 => "0000000000000000",
60057 => "0000000000000000",60058 => "0000000000000000",
60059 => "0000000000000000",60060 => "0000000000000000",
60061 => "0000000000000000",60062 => "0000000000000000",
60063 => "0000000000000000",60064 => "0000000000000000",
60065 => "0000000000000000",60066 => "0000000000000000",
60067 => "0000000000000000",60068 => "0000000000000000",
60069 => "0000000000000000",60070 => "0000000000000000",
60071 => "0000000000000000",60072 => "0000000000000000",
60073 => "0000000000000000",60074 => "0000000000000000",
60075 => "0000000000000000",60076 => "0000000000000000",
60077 => "0000000000000000",60078 => "0000000000000000",
60079 => "0000000000000000",60080 => "0000000000000000",
60081 => "0000000000000000",60082 => "0000000000000000",
60083 => "0000000000000000",60084 => "0000000000000000",
60085 => "0000000000000000",60086 => "0000000000000000",
60087 => "0000000000000000",60088 => "0000000000000000",
60089 => "0000000000000000",60090 => "0000000000000000",
60091 => "0000000000000000",60092 => "0000000000000000",
60093 => "0000000000000000",60094 => "0000000000000000",
60095 => "0000000000000000",60096 => "0000000000000000",
60097 => "0000000000000000",60098 => "0000000000000000",
60099 => "0000000000000000",60100 => "0000000000000000",
60101 => "0000000000000000",60102 => "0000000000000000",
60103 => "0000000000000000",60104 => "0000000000000000",
60105 => "0000000000000000",60106 => "0000000000000000",
60107 => "0000000000000000",60108 => "0000000000000000",
60109 => "0000000000000000",60110 => "0000000000000000",
60111 => "0000000000000000",60112 => "0000000000000000",
60113 => "0000000000000000",60114 => "0000000000000000",
60115 => "0000000000000000",60116 => "0000000000000000",
60117 => "0000000000000000",60118 => "0000000000000000",
60119 => "0000000000000000",60120 => "0000000000000000",
60121 => "0000000000000000",60122 => "0000000000000000",
60123 => "0000000000000000",60124 => "0000000000000000",
60125 => "0000000000000000",60126 => "0000000000000000",
60127 => "0000000000000000",60128 => "0000000000000000",
60129 => "0000000000000000",60130 => "0000000000000000",
60131 => "0000000000000000",60132 => "0000000000000000",
60133 => "0000000000000000",60134 => "0000000000000000",
60135 => "0000000000000000",60136 => "0000000000000000",
60137 => "0000000000000000",60138 => "0000000000000000",
60139 => "0000000000000000",60140 => "0000000000000000",
60141 => "0000000000000000",60142 => "0000000000000000",
60143 => "0000000000000000",60144 => "0000000000000000",
60145 => "0000000000000000",60146 => "0000000000000000",
60147 => "0000000000000000",60148 => "0000000000000000",
60149 => "0000000000000000",60150 => "0000000000000000",
60151 => "0000000000000000",60152 => "0000000000000000",
60153 => "0000000000000000",60154 => "0000000000000000",
60155 => "0000000000000000",60156 => "0000000000000000",
60157 => "0000000000000000",60158 => "0000000000000000",
60159 => "0000000000000000",60160 => "0000000000000000",
60161 => "0000000000000000",60162 => "0000000000000000",
60163 => "0000000000000000",60164 => "0000000000000000",
60165 => "0000000000000000",60166 => "0000000000000000",
60167 => "0000000000000000",60168 => "0000000000000000",
60169 => "0000000000000000",60170 => "0000000000000000",
60171 => "0000000000000000",60172 => "0000000000000000",
60173 => "0000000000000000",60174 => "0000000000000000",
60175 => "0000000000000000",60176 => "0000000000000000",
60177 => "0000000000000000",60178 => "0000000000000000",
60179 => "0000000000000000",60180 => "0000000000000000",
60181 => "0000000000000000",60182 => "0000000000000000",
60183 => "0000000000000000",60184 => "0000000000000000",
60185 => "0000000000000000",60186 => "0000000000000000",
60187 => "0000000000000000",60188 => "0000000000000000",
60189 => "0000000000000000",60190 => "0000000000000000",
60191 => "0000000000000000",60192 => "0000000000000000",
60193 => "0000000000000000",60194 => "0000000000000000",
60195 => "0000000000000000",60196 => "0000000000000000",
60197 => "0000000000000000",60198 => "0000000000000000",
60199 => "0000000000000000",60200 => "0000000000000000",
60201 => "0000000000000000",60202 => "0000000000000000",
60203 => "0000000000000000",60204 => "0000000000000000",
60205 => "0000000000000000",60206 => "0000000000000000",
60207 => "0000000000000000",60208 => "0000000000000000",
60209 => "0000000000000000",60210 => "0000000000000000",
60211 => "0000000000000000",60212 => "0000000000000000",
60213 => "0000000000000000",60214 => "0000000000000000",
60215 => "0000000000000000",60216 => "0000000000000000",
60217 => "0000000000000000",60218 => "0000000000000000",
60219 => "0000000000000000",60220 => "0000000000000000",
60221 => "0000000000000000",60222 => "0000000000000000",
60223 => "0000000000000000",60224 => "0000000000000000",
60225 => "0000000000000000",60226 => "0000000000000000",
60227 => "0000000000000000",60228 => "0000000000000000",
60229 => "0000000000000000",60230 => "0000000000000000",
60231 => "0000000000000000",60232 => "0000000000000000",
60233 => "0000000000000000",60234 => "0000000000000000",
60235 => "0000000000000000",60236 => "0000000000000000",
60237 => "0000000000000000",60238 => "0000000000000000",
60239 => "0000000000000000",60240 => "0000000000000000",
60241 => "0000000000000000",60242 => "0000000000000000",
60243 => "0000000000000000",60244 => "0000000000000000",
60245 => "0000000000000000",60246 => "0000000000000000",
60247 => "0000000000000000",60248 => "0000000000000000",
60249 => "0000000000000000",60250 => "0000000000000000",
60251 => "0000000000000000",60252 => "0000000000000000",
60253 => "0000000000000000",60254 => "0000000000000000",
60255 => "0000000000000000",60256 => "0000000000000000",
60257 => "0000000000000000",60258 => "0000000000000000",
60259 => "0000000000000000",60260 => "0000000000000000",
60261 => "0000000000000000",60262 => "0000000000000000",
60263 => "0000000000000000",60264 => "0000000000000000",
60265 => "0000000000000000",60266 => "0000000000000000",
60267 => "0000000000000000",60268 => "0000000000000000",
60269 => "0000000000000000",60270 => "0000000000000000",
60271 => "0000000000000000",60272 => "0000000000000000",
60273 => "0000000000000000",60274 => "0000000000000000",
60275 => "0000000000000000",60276 => "0000000000000000",
60277 => "0000000000000000",60278 => "0000000000000000",
60279 => "0000000000000000",60280 => "0000000000000000",
60281 => "0000000000000000",60282 => "0000000000000000",
60283 => "0000000000000000",60284 => "0000000000000000",
60285 => "0000000000000000",60286 => "0000000000000000",
60287 => "0000000000000000",60288 => "0000000000000000",
60289 => "0000000000000000",60290 => "0000000000000000",
60291 => "0000000000000000",60292 => "0000000000000000",
60293 => "0000000000000000",60294 => "0000000000000000",
60295 => "0000000000000000",60296 => "0000000000000000",
60297 => "0000000000000000",60298 => "0000000000000000",
60299 => "0000000000000000",60300 => "0000000000000000",
60301 => "0000000000000000",60302 => "0000000000000000",
60303 => "0000000000000000",60304 => "0000000000000000",
60305 => "0000000000000000",60306 => "0000000000000000",
60307 => "0000000000000000",60308 => "0000000000000000",
60309 => "0000000000000000",60310 => "0000000000000000",
60311 => "0000000000000000",60312 => "0000000000000000",
60313 => "0000000000000000",60314 => "0000000000000000",
60315 => "0000000000000000",60316 => "0000000000000000",
60317 => "0000000000000000",60318 => "0000000000000000",
60319 => "0000000000000000",60320 => "0000000000000000",
60321 => "0000000000000000",60322 => "0000000000000000",
60323 => "0000000000000000",60324 => "0000000000000000",
60325 => "0000000000000000",60326 => "0000000000000000",
60327 => "0000000000000000",60328 => "0000000000000000",
60329 => "0000000000000000",60330 => "0000000000000000",
60331 => "0000000000000000",60332 => "0000000000000000",
60333 => "0000000000000000",60334 => "0000000000000000",
60335 => "0000000000000000",60336 => "0000000000000000",
60337 => "0000000000000000",60338 => "0000000000000000",
60339 => "0000000000000000",60340 => "0000000000000000",
60341 => "0000000000000000",60342 => "0000000000000000",
60343 => "0000000000000000",60344 => "0000000000000000",
60345 => "0000000000000000",60346 => "0000000000000000",
60347 => "0000000000000000",60348 => "0000000000000000",
60349 => "0000000000000000",60350 => "0000000000000000",
60351 => "0000000000000000",60352 => "0000000000000000",
60353 => "0000000000000000",60354 => "0000000000000000",
60355 => "0000000000000000",60356 => "0000000000000000",
60357 => "0000000000000000",60358 => "0000000000000000",
60359 => "0000000000000000",60360 => "0000000000000000",
60361 => "0000000000000000",60362 => "0000000000000000",
60363 => "0000000000000000",60364 => "0000000000000000",
60365 => "0000000000000000",60366 => "0000000000000000",
60367 => "0000000000000000",60368 => "0000000000000000",
60369 => "0000000000000000",60370 => "0000000000000000",
60371 => "0000000000000000",60372 => "0000000000000000",
60373 => "0000000000000000",60374 => "0000000000000000",
60375 => "0000000000000000",60376 => "0000000000000000",
60377 => "0000000000000000",60378 => "0000000000000000",
60379 => "0000000000000000",60380 => "0000000000000000",
60381 => "0000000000000000",60382 => "0000000000000000",
60383 => "0000000000000000",60384 => "0000000000000000",
60385 => "0000000000000000",60386 => "0000000000000000",
60387 => "0000000000000000",60388 => "0000000000000000",
60389 => "0000000000000000",60390 => "0000000000000000",
60391 => "0000000000000000",60392 => "0000000000000000",
60393 => "0000000000000000",60394 => "0000000000000000",
60395 => "0000000000000000",60396 => "0000000000000000",
60397 => "0000000000000000",60398 => "0000000000000000",
60399 => "0000000000000000",60400 => "0000000000000000",
60401 => "0000000000000000",60402 => "0000000000000000",
60403 => "0000000000000000",60404 => "0000000000000000",
60405 => "0000000000000000",60406 => "0000000000000000",
60407 => "0000000000000000",60408 => "0000000000000000",
60409 => "0000000000000000",60410 => "0000000000000000",
60411 => "0000000000000000",60412 => "0000000000000000",
60413 => "0000000000000000",60414 => "0000000000000000",
60415 => "0000000000000000",60416 => "0000000000000000",
60417 => "0000000000000000",60418 => "0000000000000000",
60419 => "0000000000000000",60420 => "0000000000000000",
60421 => "0000000000000000",60422 => "0000000000000000",
60423 => "0000000000000000",60424 => "0000000000000000",
60425 => "0000000000000000",60426 => "0000000000000000",
60427 => "0000000000000000",60428 => "0000000000000000",
60429 => "0000000000000000",60430 => "0000000000000000",
60431 => "0000000000000000",60432 => "0000000000000000",
60433 => "0000000000000000",60434 => "0000000000000000",
60435 => "0000000000000000",60436 => "0000000000000000",
60437 => "0000000000000000",60438 => "0000000000000000",
60439 => "0000000000000000",60440 => "0000000000000000",
60441 => "0000000000000000",60442 => "0000000000000000",
60443 => "0000000000000000",60444 => "0000000000000000",
60445 => "0000000000000000",60446 => "0000000000000000",
60447 => "0000000000000000",60448 => "0000000000000000",
60449 => "0000000000000000",60450 => "0000000000000000",
60451 => "0000000000000000",60452 => "0000000000000000",
60453 => "0000000000000000",60454 => "0000000000000000",
60455 => "0000000000000000",60456 => "0000000000000000",
60457 => "0000000000000000",60458 => "0000000000000000",
60459 => "0000000000000000",60460 => "0000000000000000",
60461 => "0000000000000000",60462 => "0000000000000000",
60463 => "0000000000000000",60464 => "0000000000000000",
60465 => "0000000000000000",60466 => "0000000000000000",
60467 => "0000000000000000",60468 => "0000000000000000",
60469 => "0000000000000000",60470 => "0000000000000000",
60471 => "0000000000000000",60472 => "0000000000000000",
60473 => "0000000000000000",60474 => "0000000000000000",
60475 => "0000000000000000",60476 => "0000000000000000",
60477 => "0000000000000000",60478 => "0000000000000000",
60479 => "0000000000000000",60480 => "0000000000000000",
60481 => "0000000000000000",60482 => "0000000000000000",
60483 => "0000000000000000",60484 => "0000000000000000",
60485 => "0000000000000000",60486 => "0000000000000000",
60487 => "0000000000000000",60488 => "0000000000000000",
60489 => "0000000000000000",60490 => "0000000000000000",
60491 => "0000000000000000",60492 => "0000000000000000",
60493 => "0000000000000000",60494 => "0000000000000000",
60495 => "0000000000000000",60496 => "0000000000000000",
60497 => "0000000000000000",60498 => "0000000000000000",
60499 => "0000000000000000",60500 => "0000000000000000",
60501 => "0000000000000000",60502 => "0000000000000000",
60503 => "0000000000000000",60504 => "0000000000000000",
60505 => "0000000000000000",60506 => "0000000000000000",
60507 => "0000000000000000",60508 => "0000000000000000",
60509 => "0000000000000000",60510 => "0000000000000000",
60511 => "0000000000000000",60512 => "0000000000000000",
60513 => "0000000000000000",60514 => "0000000000000000",
60515 => "0000000000000000",60516 => "0000000000000000",
60517 => "0000000000000000",60518 => "0000000000000000",
60519 => "0000000000000000",60520 => "0000000000000000",
60521 => "0000000000000000",60522 => "0000000000000000",
60523 => "0000000000000000",60524 => "0000000000000000",
60525 => "0000000000000000",60526 => "0000000000000000",
60527 => "0000000000000000",60528 => "0000000000000000",
60529 => "0000000000000000",60530 => "0000000000000000",
60531 => "0000000000000000",60532 => "0000000000000000",
60533 => "0000000000000000",60534 => "0000000000000000",
60535 => "0000000000000000",60536 => "0000000000000000",
60537 => "0000000000000000",60538 => "0000000000000000",
60539 => "0000000000000000",60540 => "0000000000000000",
60541 => "0000000000000000",60542 => "0000000000000000",
60543 => "0000000000000000",60544 => "0000000000000000",
60545 => "0000000000000000",60546 => "0000000000000000",
60547 => "0000000000000000",60548 => "0000000000000000",
60549 => "0000000000000000",60550 => "0000000000000000",
60551 => "0000000000000000",60552 => "0000000000000000",
60553 => "0000000000000000",60554 => "0000000000000000",
60555 => "0000000000000000",60556 => "0000000000000000",
60557 => "0000000000000000",60558 => "0000000000000000",
60559 => "0000000000000000",60560 => "0000000000000000",
60561 => "0000000000000000",60562 => "0000000000000000",
60563 => "0000000000000000",60564 => "0000000000000000",
60565 => "0000000000000000",60566 => "0000000000000000",
60567 => "0000000000000000",60568 => "0000000000000000",
60569 => "0000000000000000",60570 => "0000000000000000",
60571 => "0000000000000000",60572 => "0000000000000000",
60573 => "0000000000000000",60574 => "0000000000000000",
60575 => "0000000000000000",60576 => "0000000000000000",
60577 => "0000000000000000",60578 => "0000000000000000",
60579 => "0000000000000000",60580 => "0000000000000000",
60581 => "0000000000000000",60582 => "0000000000000000",
60583 => "0000000000000000",60584 => "0000000000000000",
60585 => "0000000000000000",60586 => "0000000000000000",
60587 => "0000000000000000",60588 => "0000000000000000",
60589 => "0000000000000000",60590 => "0000000000000000",
60591 => "0000000000000000",60592 => "0000000000000000",
60593 => "0000000000000000",60594 => "0000000000000000",
60595 => "0000000000000000",60596 => "0000000000000000",
60597 => "0000000000000000",60598 => "0000000000000000",
60599 => "0000000000000000",60600 => "0000000000000000",
60601 => "0000000000000000",60602 => "0000000000000000",
60603 => "0000000000000000",60604 => "0000000000000000",
60605 => "0000000000000000",60606 => "0000000000000000",
60607 => "0000000000000000",60608 => "0000000000000000",
60609 => "0000000000000000",60610 => "0000000000000000",
60611 => "0000000000000000",60612 => "0000000000000000",
60613 => "0000000000000000",60614 => "0000000000000000",
60615 => "0000000000000000",60616 => "0000000000000000",
60617 => "0000000000000000",60618 => "0000000000000000",
60619 => "0000000000000000",60620 => "0000000000000000",
60621 => "0000000000000000",60622 => "0000000000000000",
60623 => "0000000000000000",60624 => "0000000000000000",
60625 => "0000000000000000",60626 => "0000000000000000",
60627 => "0000000000000000",60628 => "0000000000000000",
60629 => "0000000000000000",60630 => "0000000000000000",
60631 => "0000000000000000",60632 => "0000000000000000",
60633 => "0000000000000000",60634 => "0000000000000000",
60635 => "0000000000000000",60636 => "0000000000000000",
60637 => "0000000000000000",60638 => "0000000000000000",
60639 => "0000000000000000",60640 => "0000000000000000",
60641 => "0000000000000000",60642 => "0000000000000000",
60643 => "0000000000000000",60644 => "0000000000000000",
60645 => "0000000000000000",60646 => "0000000000000000",
60647 => "0000000000000000",60648 => "0000000000000000",
60649 => "0000000000000000",60650 => "0000000000000000",
60651 => "0000000000000000",60652 => "0000000000000000",
60653 => "0000000000000000",60654 => "0000000000000000",
60655 => "0000000000000000",60656 => "0000000000000000",
60657 => "0000000000000000",60658 => "0000000000000000",
60659 => "0000000000000000",60660 => "0000000000000000",
60661 => "0000000000000000",60662 => "0000000000000000",
60663 => "0000000000000000",60664 => "0000000000000000",
60665 => "0000000000000000",60666 => "0000000000000000",
60667 => "0000000000000000",60668 => "0000000000000000",
60669 => "0000000000000000",60670 => "0000000000000000",
60671 => "0000000000000000",60672 => "0000000000000000",
60673 => "0000000000000000",60674 => "0000000000000000",
60675 => "0000000000000000",60676 => "0000000000000000",
60677 => "0000000000000000",60678 => "0000000000000000",
60679 => "0000000000000000",60680 => "0000000000000000",
60681 => "0000000000000000",60682 => "0000000000000000",
60683 => "0000000000000000",60684 => "0000000000000000",
60685 => "0000000000000000",60686 => "0000000000000000",
60687 => "0000000000000000",60688 => "0000000000000000",
60689 => "0000000000000000",60690 => "0000000000000000",
60691 => "0000000000000000",60692 => "0000000000000000",
60693 => "0000000000000000",60694 => "0000000000000000",
60695 => "0000000000000000",60696 => "0000000000000000",
60697 => "0000000000000000",60698 => "0000000000000000",
60699 => "0000000000000000",60700 => "0000000000000000",
60701 => "0000000000000000",60702 => "0000000000000000",
60703 => "0000000000000000",60704 => "0000000000000000",
60705 => "0000000000000000",60706 => "0000000000000000",
60707 => "0000000000000000",60708 => "0000000000000000",
60709 => "0000000000000000",60710 => "0000000000000000",
60711 => "0000000000000000",60712 => "0000000000000000",
60713 => "0000000000000000",60714 => "0000000000000000",
60715 => "0000000000000000",60716 => "0000000000000000",
60717 => "0000000000000000",60718 => "0000000000000000",
60719 => "0000000000000000",60720 => "0000000000000000",
60721 => "0000000000000000",60722 => "0000000000000000",
60723 => "0000000000000000",60724 => "0000000000000000",
60725 => "0000000000000000",60726 => "0000000000000000",
60727 => "0000000000000000",60728 => "0000000000000000",
60729 => "0000000000000000",60730 => "0000000000000000",
60731 => "0000000000000000",60732 => "0000000000000000",
60733 => "0000000000000000",60734 => "0000000000000000",
60735 => "0000000000000000",60736 => "0000000000000000",
60737 => "0000000000000000",60738 => "0000000000000000",
60739 => "0000000000000000",60740 => "0000000000000000",
60741 => "0000000000000000",60742 => "0000000000000000",
60743 => "0000000000000000",60744 => "0000000000000000",
60745 => "0000000000000000",60746 => "0000000000000000",
60747 => "0000000000000000",60748 => "0000000000000000",
60749 => "0000000000000000",60750 => "0000000000000000",
60751 => "0000000000000000",60752 => "0000000000000000",
60753 => "0000000000000000",60754 => "0000000000000000",
60755 => "0000000000000000",60756 => "0000000000000000",
60757 => "0000000000000000",60758 => "0000000000000000",
60759 => "0000000000000000",60760 => "0000000000000000",
60761 => "0000000000000000",60762 => "0000000000000000",
60763 => "0000000000000000",60764 => "0000000000000000",
60765 => "0000000000000000",60766 => "0000000000000000",
60767 => "0000000000000000",60768 => "0000000000000000",
60769 => "0000000000000000",60770 => "0000000000000000",
60771 => "0000000000000000",60772 => "0000000000000000",
60773 => "0000000000000000",60774 => "0000000000000000",
60775 => "0000000000000000",60776 => "0000000000000000",
60777 => "0000000000000000",60778 => "0000000000000000",
60779 => "0000000000000000",60780 => "0000000000000000",
60781 => "0000000000000000",60782 => "0000000000000000",
60783 => "0000000000000000",60784 => "0000000000000000",
60785 => "0000000000000000",60786 => "0000000000000000",
60787 => "0000000000000000",60788 => "0000000000000000",
60789 => "0000000000000000",60790 => "0000000000000000",
60791 => "0000000000000000",60792 => "0000000000000000",
60793 => "0000000000000000",60794 => "0000000000000000",
60795 => "0000000000000000",60796 => "0000000000000000",
60797 => "0000000000000000",60798 => "0000000000000000",
60799 => "0000000000000000",60800 => "0000000000000000",
60801 => "0000000000000000",60802 => "0000000000000000",
60803 => "0000000000000000",60804 => "0000000000000000",
60805 => "0000000000000000",60806 => "0000000000000000",
60807 => "0000000000000000",60808 => "0000000000000000",
60809 => "0000000000000000",60810 => "0000000000000000",
60811 => "0000000000000000",60812 => "0000000000000000",
60813 => "0000000000000000",60814 => "0000000000000000",
60815 => "0000000000000000",60816 => "0000000000000000",
60817 => "0000000000000000",60818 => "0000000000000000",
60819 => "0000000000000000",60820 => "0000000000000000",
60821 => "0000000000000000",60822 => "0000000000000000",
60823 => "0000000000000000",60824 => "0000000000000000",
60825 => "0000000000000000",60826 => "0000000000000000",
60827 => "0000000000000000",60828 => "0000000000000000",
60829 => "0000000000000000",60830 => "0000000000000000",
60831 => "0000000000000000",60832 => "0000000000000000",
60833 => "0000000000000000",60834 => "0000000000000000",
60835 => "0000000000000000",60836 => "0000000000000000",
60837 => "0000000000000000",60838 => "0000000000000000",
60839 => "0000000000000000",60840 => "0000000000000000",
60841 => "0000000000000000",60842 => "0000000000000000",
60843 => "0000000000000000",60844 => "0000000000000000",
60845 => "0000000000000000",60846 => "0000000000000000",
60847 => "0000000000000000",60848 => "0000000000000000",
60849 => "0000000000000000",60850 => "0000000000000000",
60851 => "0000000000000000",60852 => "0000000000000000",
60853 => "0000000000000000",60854 => "0000000000000000",
60855 => "0000000000000000",60856 => "0000000000000000",
60857 => "0000000000000000",60858 => "0000000000000000",
60859 => "0000000000000000",60860 => "0000000000000000",
60861 => "0000000000000000",60862 => "0000000000000000",
60863 => "0000000000000000",60864 => "0000000000000000",
60865 => "0000000000000000",60866 => "0000000000000000",
60867 => "0000000000000000",60868 => "0000000000000000",
60869 => "0000000000000000",60870 => "0000000000000000",
60871 => "0000000000000000",60872 => "0000000000000000",
60873 => "0000000000000000",60874 => "0000000000000000",
60875 => "0000000000000000",60876 => "0000000000000000",
60877 => "0000000000000000",60878 => "0000000000000000",
60879 => "0000000000000000",60880 => "0000000000000000",
60881 => "0000000000000000",60882 => "0000000000000000",
60883 => "0000000000000000",60884 => "0000000000000000",
60885 => "0000000000000000",60886 => "0000000000000000",
60887 => "0000000000000000",60888 => "0000000000000000",
60889 => "0000000000000000",60890 => "0000000000000000",
60891 => "0000000000000000",60892 => "0000000000000000",
60893 => "0000000000000000",60894 => "0000000000000000",
60895 => "0000000000000000",60896 => "0000000000000000",
60897 => "0000000000000000",60898 => "0000000000000000",
60899 => "0000000000000000",60900 => "0000000000000000",
60901 => "0000000000000000",60902 => "0000000000000000",
60903 => "0000000000000000",60904 => "0000000000000000",
60905 => "0000000000000000",60906 => "0000000000000000",
60907 => "0000000000000000",60908 => "0000000000000000",
60909 => "0000000000000000",60910 => "0000000000000000",
60911 => "0000000000000000",60912 => "0000000000000000",
60913 => "0000000000000000",60914 => "0000000000000000",
60915 => "0000000000000000",60916 => "0000000000000000",
60917 => "0000000000000000",60918 => "0000000000000000",
60919 => "0000000000000000",60920 => "0000000000000000",
60921 => "0000000000000000",60922 => "0000000000000000",
60923 => "0000000000000000",60924 => "0000000000000000",
60925 => "0000000000000000",60926 => "0000000000000000",
60927 => "0000000000000000",60928 => "0000000000000000",
60929 => "0000000000000000",60930 => "0000000000000000",
60931 => "0000000000000000",60932 => "0000000000000000",
60933 => "0000000000000000",60934 => "0000000000000000",
60935 => "0000000000000000",60936 => "0000000000000000",
60937 => "0000000000000000",60938 => "0000000000000000",
60939 => "0000000000000000",60940 => "0000000000000000",
60941 => "0000000000000000",60942 => "0000000000000000",
60943 => "0000000000000000",60944 => "0000000000000000",
60945 => "0000000000000000",60946 => "0000000000000000",
60947 => "0000000000000000",60948 => "0000000000000000",
60949 => "0000000000000000",60950 => "0000000000000000",
60951 => "0000000000000000",60952 => "0000000000000000",
60953 => "0000000000000000",60954 => "0000000000000000",
60955 => "0000000000000000",60956 => "0000000000000000",
60957 => "0000000000000000",60958 => "0000000000000000",
60959 => "0000000000000000",60960 => "0000000000000000",
60961 => "0000000000000000",60962 => "0000000000000000",
60963 => "0000000000000000",60964 => "0000000000000000",
60965 => "0000000000000000",60966 => "0000000000000000",
60967 => "0000000000000000",60968 => "0000000000000000",
60969 => "0000000000000000",60970 => "0000000000000000",
60971 => "0000000000000000",60972 => "0000000000000000",
60973 => "0000000000000000",60974 => "0000000000000000",
60975 => "0000000000000000",60976 => "0000000000000000",
60977 => "0000000000000000",60978 => "0000000000000000",
60979 => "0000000000000000",60980 => "0000000000000000",
60981 => "0000000000000000",60982 => "0000000000000000",
60983 => "0000000000000000",60984 => "0000000000000000",
60985 => "0000000000000000",60986 => "0000000000000000",
60987 => "0000000000000000",60988 => "0000000000000000",
60989 => "0000000000000000",60990 => "0000000000000000",
60991 => "0000000000000000",60992 => "0000000000000000",
60993 => "0000000000000000",60994 => "0000000000000000",
60995 => "0000000000000000",60996 => "0000000000000000",
60997 => "0000000000000000",60998 => "0000000000000000",
60999 => "0000000000000000",61000 => "0000000000000000",
61001 => "0000000000000000",61002 => "0000000000000000",
61003 => "0000000000000000",61004 => "0000000000000000",
61005 => "0000000000000000",61006 => "0000000000000000",
61007 => "0000000000000000",61008 => "0000000000000000",
61009 => "0000000000000000",61010 => "0000000000000000",
61011 => "0000000000000000",61012 => "0000000000000000",
61013 => "0000000000000000",61014 => "0000000000000000",
61015 => "0000000000000000",61016 => "0000000000000000",
61017 => "0000000000000000",61018 => "0000000000000000",
61019 => "0000000000000000",61020 => "0000000000000000",
61021 => "0000000000000000",61022 => "0000000000000000",
61023 => "0000000000000000",61024 => "0000000000000000",
61025 => "0000000000000000",61026 => "0000000000000000",
61027 => "0000000000000000",61028 => "0000000000000000",
61029 => "0000000000000000",61030 => "0000000000000000",
61031 => "0000000000000000",61032 => "0000000000000000",
61033 => "0000000000000000",61034 => "0000000000000000",
61035 => "0000000000000000",61036 => "0000000000000000",
61037 => "0000000000000000",61038 => "0000000000000000",
61039 => "0000000000000000",61040 => "0000000000000000",
61041 => "0000000000000000",61042 => "0000000000000000",
61043 => "0000000000000000",61044 => "0000000000000000",
61045 => "0000000000000000",61046 => "0000000000000000",
61047 => "0000000000000000",61048 => "0000000000000000",
61049 => "0000000000000000",61050 => "0000000000000000",
61051 => "0000000000000000",61052 => "0000000000000000",
61053 => "0000000000000000",61054 => "0000000000000000",
61055 => "0000000000000000",61056 => "0000000000000000",
61057 => "0000000000000000",61058 => "0000000000000000",
61059 => "0000000000000000",61060 => "0000000000000000",
61061 => "0000000000000000",61062 => "0000000000000000",
61063 => "0000000000000000",61064 => "0000000000000000",
61065 => "0000000000000000",61066 => "0000000000000000",
61067 => "0000000000000000",61068 => "0000000000000000",
61069 => "0000000000000000",61070 => "0000000000000000",
61071 => "0000000000000000",61072 => "0000000000000000",
61073 => "0000000000000000",61074 => "0000000000000000",
61075 => "0000000000000000",61076 => "0000000000000000",
61077 => "0000000000000000",61078 => "0000000000000000",
61079 => "0000000000000000",61080 => "0000000000000000",
61081 => "0000000000000000",61082 => "0000000000000000",
61083 => "0000000000000000",61084 => "0000000000000000",
61085 => "0000000000000000",61086 => "0000000000000000",
61087 => "0000000000000000",61088 => "0000000000000000",
61089 => "0000000000000000",61090 => "0000000000000000",
61091 => "0000000000000000",61092 => "0000000000000000",
61093 => "0000000000000000",61094 => "0000000000000000",
61095 => "0000000000000000",61096 => "0000000000000000",
61097 => "0000000000000000",61098 => "0000000000000000",
61099 => "0000000000000000",61100 => "0000000000000000",
61101 => "0000000000000000",61102 => "0000000000000000",
61103 => "0000000000000000",61104 => "0000000000000000",
61105 => "0000000000000000",61106 => "0000000000000000",
61107 => "0000000000000000",61108 => "0000000000000000",
61109 => "0000000000000000",61110 => "0000000000000000",
61111 => "0000000000000000",61112 => "0000000000000000",
61113 => "0000000000000000",61114 => "0000000000000000",
61115 => "0000000000000000",61116 => "0000000000000000",
61117 => "0000000000000000",61118 => "0000000000000000",
61119 => "0000000000000000",61120 => "0000000000000000",
61121 => "0000000000000000",61122 => "0000000000000000",
61123 => "0000000000000000",61124 => "0000000000000000",
61125 => "0000000000000000",61126 => "0000000000000000",
61127 => "0000000000000000",61128 => "0000000000000000",
61129 => "0000000000000000",61130 => "0000000000000000",
61131 => "0000000000000000",61132 => "0000000000000000",
61133 => "0000000000000000",61134 => "0000000000000000",
61135 => "0000000000000000",61136 => "0000000000000000",
61137 => "0000000000000000",61138 => "0000000000000000",
61139 => "0000000000000000",61140 => "0000000000000000",
61141 => "0000000000000000",61142 => "0000000000000000",
61143 => "0000000000000000",61144 => "0000000000000000",
61145 => "0000000000000000",61146 => "0000000000000000",
61147 => "0000000000000000",61148 => "0000000000000000",
61149 => "0000000000000000",61150 => "0000000000000000",
61151 => "0000000000000000",61152 => "0000000000000000",
61153 => "0000000000000000",61154 => "0000000000000000",
61155 => "0000000000000000",61156 => "0000000000000000",
61157 => "0000000000000000",61158 => "0000000000000000",
61159 => "0000000000000000",61160 => "0000000000000000",
61161 => "0000000000000000",61162 => "0000000000000000",
61163 => "0000000000000000",61164 => "0000000000000000",
61165 => "0000000000000000",61166 => "0000000000000000",
61167 => "0000000000000000",61168 => "0000000000000000",
61169 => "0000000000000000",61170 => "0000000000000000",
61171 => "0000000000000000",61172 => "0000000000000000",
61173 => "0000000000000000",61174 => "0000000000000000",
61175 => "0000000000000000",61176 => "0000000000000000",
61177 => "0000000000000000",61178 => "0000000000000000",
61179 => "0000000000000000",61180 => "0000000000000000",
61181 => "0000000000000000",61182 => "0000000000000000",
61183 => "0000000000000000",61184 => "0000000000000000",
61185 => "0000000000000000",61186 => "0000000000000000",
61187 => "0000000000000000",61188 => "0000000000000000",
61189 => "0000000000000000",61190 => "0000000000000000",
61191 => "0000000000000000",61192 => "0000000000000000",
61193 => "0000000000000000",61194 => "0000000000000000",
61195 => "0000000000000000",61196 => "0000000000000000",
61197 => "0000000000000000",61198 => "0000000000000000",
61199 => "0000000000000000",61200 => "0000000000000000",
61201 => "0000000000000000",61202 => "0000000000000000",
61203 => "0000000000000000",61204 => "0000000000000000",
61205 => "0000000000000000",61206 => "0000000000000000",
61207 => "0000000000000000",61208 => "0000000000000000",
61209 => "0000000000000000",61210 => "0000000000000000",
61211 => "0000000000000000",61212 => "0000000000000000",
61213 => "0000000000000000",61214 => "0000000000000000",
61215 => "0000000000000000",61216 => "0000000000000000",
61217 => "0000000000000000",61218 => "0000000000000000",
61219 => "0000000000000000",61220 => "0000000000000000",
61221 => "0000000000000000",61222 => "0000000000000000",
61223 => "0000000000000000",61224 => "0000000000000000",
61225 => "0000000000000000",61226 => "0000000000000000",
61227 => "0000000000000000",61228 => "0000000000000000",
61229 => "0000000000000000",61230 => "0000000000000000",
61231 => "0000000000000000",61232 => "0000000000000000",
61233 => "0000000000000000",61234 => "0000000000000000",
61235 => "0000000000000000",61236 => "0000000000000000",
61237 => "0000000000000000",61238 => "0000000000000000",
61239 => "0000000000000000",61240 => "0000000000000000",
61241 => "0000000000000000",61242 => "0000000000000000",
61243 => "0000000000000000",61244 => "0000000000000000",
61245 => "0000000000000000",61246 => "0000000000000000",
61247 => "0000000000000000",61248 => "0000000000000000",
61249 => "0000000000000000",61250 => "0000000000000000",
61251 => "0000000000000000",61252 => "0000000000000000",
61253 => "0000000000000000",61254 => "0000000000000000",
61255 => "0000000000000000",61256 => "0000000000000000",
61257 => "0000000000000000",61258 => "0000000000000000",
61259 => "0000000000000000",61260 => "0000000000000000",
61261 => "0000000000000000",61262 => "0000000000000000",
61263 => "0000000000000000",61264 => "0000000000000000",
61265 => "0000000000000000",61266 => "0000000000000000",
61267 => "0000000000000000",61268 => "0000000000000000",
61269 => "0000000000000000",61270 => "0000000000000000",
61271 => "0000000000000000",61272 => "0000000000000000",
61273 => "0000000000000000",61274 => "0000000000000000",
61275 => "0000000000000000",61276 => "0000000000000000",
61277 => "0000000000000000",61278 => "0000000000000000",
61279 => "0000000000000000",61280 => "0000000000000000",
61281 => "0000000000000000",61282 => "0000000000000000",
61283 => "0000000000000000",61284 => "0000000000000000",
61285 => "0000000000000000",61286 => "0000000000000000",
61287 => "0000000000000000",61288 => "0000000000000000",
61289 => "0000000000000000",61290 => "0000000000000000",
61291 => "0000000000000000",61292 => "0000000000000000",
61293 => "0000000000000000",61294 => "0000000000000000",
61295 => "0000000000000000",61296 => "0000000000000000",
61297 => "0000000000000000",61298 => "0000000000000000",
61299 => "0000000000000000",61300 => "0000000000000000",
61301 => "0000000000000000",61302 => "0000000000000000",
61303 => "0000000000000000",61304 => "0000000000000000",
61305 => "0000000000000000",61306 => "0000000000000000",
61307 => "0000000000000000",61308 => "0000000000000000",
61309 => "0000000000000000",61310 => "0000000000000000",
61311 => "0000000000000000",61312 => "0000000000000000",
61313 => "0000000000000000",61314 => "0000000000000000",
61315 => "0000000000000000",61316 => "0000000000000000",
61317 => "0000000000000000",61318 => "0000000000000000",
61319 => "0000000000000000",61320 => "0000000000000000",
61321 => "0000000000000000",61322 => "0000000000000000",
61323 => "0000000000000000",61324 => "0000000000000000",
61325 => "0000000000000000",61326 => "0000000000000000",
61327 => "0000000000000000",61328 => "0000000000000000",
61329 => "0000000000000000",61330 => "0000000000000000",
61331 => "0000000000000000",61332 => "0000000000000000",
61333 => "0000000000000000",61334 => "0000000000000000",
61335 => "0000000000000000",61336 => "0000000000000000",
61337 => "0000000000000000",61338 => "0000000000000000",
61339 => "0000000000000000",61340 => "0000000000000000",
61341 => "0000000000000000",61342 => "0000000000000000",
61343 => "0000000000000000",61344 => "0000000000000000",
61345 => "0000000000000000",61346 => "0000000000000000",
61347 => "0000000000000000",61348 => "0000000000000000",
61349 => "0000000000000000",61350 => "0000000000000000",
61351 => "0000000000000000",61352 => "0000000000000000",
61353 => "0000000000000000",61354 => "0000000000000000",
61355 => "0000000000000000",61356 => "0000000000000000",
61357 => "0000000000000000",61358 => "0000000000000000",
61359 => "0000000000000000",61360 => "0000000000000000",
61361 => "0000000000000000",61362 => "0000000000000000",
61363 => "0000000000000000",61364 => "0000000000000000",
61365 => "0000000000000000",61366 => "0000000000000000",
61367 => "0000000000000000",61368 => "0000000000000000",
61369 => "0000000000000000",61370 => "0000000000000000",
61371 => "0000000000000000",61372 => "0000000000000000",
61373 => "0000000000000000",61374 => "0000000000000000",
61375 => "0000000000000000",61376 => "0000000000000000",
61377 => "0000000000000000",61378 => "0000000000000000",
61379 => "0000000000000000",61380 => "0000000000000000",
61381 => "0000000000000000",61382 => "0000000000000000",
61383 => "0000000000000000",61384 => "0000000000000000",
61385 => "0000000000000000",61386 => "0000000000000000",
61387 => "0000000000000000",61388 => "0000000000000000",
61389 => "0000000000000000",61390 => "0000000000000000",
61391 => "0000000000000000",61392 => "0000000000000000",
61393 => "0000000000000000",61394 => "0000000000000000",
61395 => "0000000000000000",61396 => "0000000000000000",
61397 => "0000000000000000",61398 => "0000000000000000",
61399 => "0000000000000000",61400 => "0000000000000000",
61401 => "0000000000000000",61402 => "0000000000000000",
61403 => "0000000000000000",61404 => "0000000000000000",
61405 => "0000000000000000",61406 => "0000000000000000",
61407 => "0000000000000000",61408 => "0000000000000000",
61409 => "0000000000000000",61410 => "0000000000000000",
61411 => "0000000000000000",61412 => "0000000000000000",
61413 => "0000000000000000",61414 => "0000000000000000",
61415 => "0000000000000000",61416 => "0000000000000000",
61417 => "0000000000000000",61418 => "0000000000000000",
61419 => "0000000000000000",61420 => "0000000000000000",
61421 => "0000000000000000",61422 => "0000000000000000",
61423 => "0000000000000000",61424 => "0000000000000000",
61425 => "0000000000000000",61426 => "0000000000000000",
61427 => "0000000000000000",61428 => "0000000000000000",
61429 => "0000000000000000",61430 => "0000000000000000",
61431 => "0000000000000000",61432 => "0000000000000000",
61433 => "0000000000000000",61434 => "0000000000000000",
61435 => "0000000000000000",61436 => "0000000000000000",
61437 => "0000000000000000",61438 => "0000000000000000",
61439 => "0000000000000000",61440 => "0000000000000000",
61441 => "0000000000000000",61442 => "0000000000000000",
61443 => "0000000000000000",61444 => "0000000000000000",
61445 => "0000000000000000",61446 => "0000000000000000",
61447 => "0000000000000000",61448 => "0000000000000000",
61449 => "0000000000000000",61450 => "0000000000000000",
61451 => "0000000000000000",61452 => "0000000000000000",
61453 => "0000000000000000",61454 => "0000000000000000",
61455 => "0000000000000000",61456 => "0000000000000000",
61457 => "0000000000000000",61458 => "0000000000000000",
61459 => "0000000000000000",61460 => "0000000000000000",
61461 => "0000000000000000",61462 => "0000000000000000",
61463 => "0000000000000000",61464 => "0000000000000000",
61465 => "0000000000000000",61466 => "0000000000000000",
61467 => "0000000000000000",61468 => "0000000000000000",
61469 => "0000000000000000",61470 => "0000000000000000",
61471 => "0000000000000000",61472 => "0000000000000000",
61473 => "0000000000000000",61474 => "0000000000000000",
61475 => "0000000000000000",61476 => "0000000000000000",
61477 => "0000000000000000",61478 => "0000000000000000",
61479 => "0000000000000000",61480 => "0000000000000000",
61481 => "0000000000000000",61482 => "0000000000000000",
61483 => "0000000000000000",61484 => "0000000000000000",
61485 => "0000000000000000",61486 => "0000000000000000",
61487 => "0000000000000000",61488 => "0000000000000000",
61489 => "0000000000000000",61490 => "0000000000000000",
61491 => "0000000000000000",61492 => "0000000000000000",
61493 => "0000000000000000",61494 => "0000000000000000",
61495 => "0000000000000000",61496 => "0000000000000000",
61497 => "0000000000000000",61498 => "0000000000000000",
61499 => "0000000000000000",61500 => "0000000000000000",
61501 => "0000000000000000",61502 => "0000000000000000",
61503 => "0000000000000000",61504 => "0000000000000000",
61505 => "0000000000000000",61506 => "0000000000000000",
61507 => "0000000000000000",61508 => "0000000000000000",
61509 => "0000000000000000",61510 => "0000000000000000",
61511 => "0000000000000000",61512 => "0000000000000000",
61513 => "0000000000000000",61514 => "0000000000000000",
61515 => "0000000000000000",61516 => "0000000000000000",
61517 => "0000000000000000",61518 => "0000000000000000",
61519 => "0000000000000000",61520 => "0000000000000000",
61521 => "0000000000000000",61522 => "0000000000000000",
61523 => "0000000000000000",61524 => "0000000000000000",
61525 => "0000000000000000",61526 => "0000000000000000",
61527 => "0000000000000000",61528 => "0000000000000000",
61529 => "0000000000000000",61530 => "0000000000000000",
61531 => "0000000000000000",61532 => "0000000000000000",
61533 => "0000000000000000",61534 => "0000000000000000",
61535 => "0000000000000000",61536 => "0000000000000000",
61537 => "0000000000000000",61538 => "0000000000000000",
61539 => "0000000000000000",61540 => "0000000000000000",
61541 => "0000000000000000",61542 => "0000000000000000",
61543 => "0000000000000000",61544 => "0000000000000000",
61545 => "0000000000000000",61546 => "0000000000000000",
61547 => "0000000000000000",61548 => "0000000000000000",
61549 => "0000000000000000",61550 => "0000000000000000",
61551 => "0000000000000000",61552 => "0000000000000000",
61553 => "0000000000000000",61554 => "0000000000000000",
61555 => "0000000000000000",61556 => "0000000000000000",
61557 => "0000000000000000",61558 => "0000000000000000",
61559 => "0000000000000000",61560 => "0000000000000000",
61561 => "0000000000000000",61562 => "0000000000000000",
61563 => "0000000000000000",61564 => "0000000000000000",
61565 => "0000000000000000",61566 => "0000000000000000",
61567 => "0000000000000000",61568 => "0000000000000000",
61569 => "0000000000000000",61570 => "0000000000000000",
61571 => "0000000000000000",61572 => "0000000000000000",
61573 => "0000000000000000",61574 => "0000000000000000",
61575 => "0000000000000000",61576 => "0000000000000000",
61577 => "0000000000000000",61578 => "0000000000000000",
61579 => "0000000000000000",61580 => "0000000000000000",
61581 => "0000000000000000",61582 => "0000000000000000",
61583 => "0000000000000000",61584 => "0000000000000000",
61585 => "0000000000000000",61586 => "0000000000000000",
61587 => "0000000000000000",61588 => "0000000000000000",
61589 => "0000000000000000",61590 => "0000000000000000",
61591 => "0000000000000000",61592 => "0000000000000000",
61593 => "0000000000000000",61594 => "0000000000000000",
61595 => "0000000000000000",61596 => "0000000000000000",
61597 => "0000000000000000",61598 => "0000000000000000",
61599 => "0000000000000000",61600 => "0000000000000000",
61601 => "0000000000000000",61602 => "0000000000000000",
61603 => "0000000000000000",61604 => "0000000000000000",
61605 => "0000000000000000",61606 => "0000000000000000",
61607 => "0000000000000000",61608 => "0000000000000000",
61609 => "0000000000000000",61610 => "0000000000000000",
61611 => "0000000000000000",61612 => "0000000000000000",
61613 => "0000000000000000",61614 => "0000000000000000",
61615 => "0000000000000000",61616 => "0000000000000000",
61617 => "0000000000000000",61618 => "0000000000000000",
61619 => "0000000000000000",61620 => "0000000000000000",
61621 => "0000000000000000",61622 => "0000000000000000",
61623 => "0000000000000000",61624 => "0000000000000000",
61625 => "0000000000000000",61626 => "0000000000000000",
61627 => "0000000000000000",61628 => "0000000000000000",
61629 => "0000000000000000",61630 => "0000000000000000",
61631 => "0000000000000000",61632 => "0000000000000000",
61633 => "0000000000000000",61634 => "0000000000000000",
61635 => "0000000000000000",61636 => "0000000000000000",
61637 => "0000000000000000",61638 => "0000000000000000",
61639 => "0000000000000000",61640 => "0000000000000000",
61641 => "0000000000000000",61642 => "0000000000000000",
61643 => "0000000000000000",61644 => "0000000000000000",
61645 => "0000000000000000",61646 => "0000000000000000",
61647 => "0000000000000000",61648 => "0000000000000000",
61649 => "0000000000000000",61650 => "0000000000000000",
61651 => "0000000000000000",61652 => "0000000000000000",
61653 => "0000000000000000",61654 => "0000000000000000",
61655 => "0000000000000000",61656 => "0000000000000000",
61657 => "0000000000000000",61658 => "0000000000000000",
61659 => "0000000000000000",61660 => "0000000000000000",
61661 => "0000000000000000",61662 => "0000000000000000",
61663 => "0000000000000000",61664 => "0000000000000000",
61665 => "0000000000000000",61666 => "0000000000000000",
61667 => "0000000000000000",61668 => "0000000000000000",
61669 => "0000000000000000",61670 => "0000000000000000",
61671 => "0000000000000000",61672 => "0000000000000000",
61673 => "0000000000000000",61674 => "0000000000000000",
61675 => "0000000000000000",61676 => "0000000000000000",
61677 => "0000000000000000",61678 => "0000000000000000",
61679 => "0000000000000000",61680 => "0000000000000000",
61681 => "0000000000000000",61682 => "0000000000000000",
61683 => "0000000000000000",61684 => "0000000000000000",
61685 => "0000000000000000",61686 => "0000000000000000",
61687 => "0000000000000000",61688 => "0000000000000000",
61689 => "0000000000000000",61690 => "0000000000000000",
61691 => "0000000000000000",61692 => "0000000000000000",
61693 => "0000000000000000",61694 => "0000000000000000",
61695 => "0000000000000000",61696 => "0000000000000000",
61697 => "0000000000000000",61698 => "0000000000000000",
61699 => "0000000000000000",61700 => "0000000000000000",
61701 => "0000000000000000",61702 => "0000000000000000",
61703 => "0000000000000000",61704 => "0000000000000000",
61705 => "0000000000000000",61706 => "0000000000000000",
61707 => "0000000000000000",61708 => "0000000000000000",
61709 => "0000000000000000",61710 => "0000000000000000",
61711 => "0000000000000000",61712 => "0000000000000000",
61713 => "0000000000000000",61714 => "0000000000000000",
61715 => "0000000000000000",61716 => "0000000000000000",
61717 => "0000000000000000",61718 => "0000000000000000",
61719 => "0000000000000000",61720 => "0000000000000000",
61721 => "0000000000000000",61722 => "0000000000000000",
61723 => "0000000000000000",61724 => "0000000000000000",
61725 => "0000000000000000",61726 => "0000000000000000",
61727 => "0000000000000000",61728 => "0000000000000000",
61729 => "0000000000000000",61730 => "0000000000000000",
61731 => "0000000000000000",61732 => "0000000000000000",
61733 => "0000000000000000",61734 => "0000000000000000",
61735 => "0000000000000000",61736 => "0000000000000000",
61737 => "0000000000000000",61738 => "0000000000000000",
61739 => "0000000000000000",61740 => "0000000000000000",
61741 => "0000000000000000",61742 => "0000000000000000",
61743 => "0000000000000000",61744 => "0000000000000000",
61745 => "0000000000000000",61746 => "0000000000000000",
61747 => "0000000000000000",61748 => "0000000000000000",
61749 => "0000000000000000",61750 => "0000000000000000",
61751 => "0000000000000000",61752 => "0000000000000000",
61753 => "0000000000000000",61754 => "0000000000000000",
61755 => "0000000000000000",61756 => "0000000000000000",
61757 => "0000000000000000",61758 => "0000000000000000",
61759 => "0000000000000000",61760 => "0000000000000000",
61761 => "0000000000000000",61762 => "0000000000000000",
61763 => "0000000000000000",61764 => "0000000000000000",
61765 => "0000000000000000",61766 => "0000000000000000",
61767 => "0000000000000000",61768 => "0000000000000000",
61769 => "0000000000000000",61770 => "0000000000000000",
61771 => "0000000000000000",61772 => "0000000000000000",
61773 => "0000000000000000",61774 => "0000000000000000",
61775 => "0000000000000000",61776 => "0000000000000000",
61777 => "0000000000000000",61778 => "0000000000000000",
61779 => "0000000000000000",61780 => "0000000000000000",
61781 => "0000000000000000",61782 => "0000000000000000",
61783 => "0000000000000000",61784 => "0000000000000000",
61785 => "0000000000000000",61786 => "0000000000000000",
61787 => "0000000000000000",61788 => "0000000000000000",
61789 => "0000000000000000",61790 => "0000000000000000",
61791 => "0000000000000000",61792 => "0000000000000000",
61793 => "0000000000000000",61794 => "0000000000000000",
61795 => "0000000000000000",61796 => "0000000000000000",
61797 => "0000000000000000",61798 => "0000000000000000",
61799 => "0000000000000000",61800 => "0000000000000000",
61801 => "0000000000000000",61802 => "0000000000000000",
61803 => "0000000000000000",61804 => "0000000000000000",
61805 => "0000000000000000",61806 => "0000000000000000",
61807 => "0000000000000000",61808 => "0000000000000000",
61809 => "0000000000000000",61810 => "0000000000000000",
61811 => "0000000000000000",61812 => "0000000000000000",
61813 => "0000000000000000",61814 => "0000000000000000",
61815 => "0000000000000000",61816 => "0000000000000000",
61817 => "0000000000000000",61818 => "0000000000000000",
61819 => "0000000000000000",61820 => "0000000000000000",
61821 => "0000000000000000",61822 => "0000000000000000",
61823 => "0000000000000000",61824 => "0000000000000000",
61825 => "0000000000000000",61826 => "0000000000000000",
61827 => "0000000000000000",61828 => "0000000000000000",
61829 => "0000000000000000",61830 => "0000000000000000",
61831 => "0000000000000000",61832 => "0000000000000000",
61833 => "0000000000000000",61834 => "0000000000000000",
61835 => "0000000000000000",61836 => "0000000000000000",
61837 => "0000000000000000",61838 => "0000000000000000",
61839 => "0000000000000000",61840 => "0000000000000000",
61841 => "0000000000000000",61842 => "0000000000000000",
61843 => "0000000000000000",61844 => "0000000000000000",
61845 => "0000000000000000",61846 => "0000000000000000",
61847 => "0000000000000000",61848 => "0000000000000000",
61849 => "0000000000000000",61850 => "0000000000000000",
61851 => "0000000000000000",61852 => "0000000000000000",
61853 => "0000000000000000",61854 => "0000000000000000",
61855 => "0000000000000000",61856 => "0000000000000000",
61857 => "0000000000000000",61858 => "0000000000000000",
61859 => "0000000000000000",61860 => "0000000000000000",
61861 => "0000000000000000",61862 => "0000000000000000",
61863 => "0000000000000000",61864 => "0000000000000000",
61865 => "0000000000000000",61866 => "0000000000000000",
61867 => "0000000000000000",61868 => "0000000000000000",
61869 => "0000000000000000",61870 => "0000000000000000",
61871 => "0000000000000000",61872 => "0000000000000000",
61873 => "0000000000000000",61874 => "0000000000000000",
61875 => "0000000000000000",61876 => "0000000000000000",
61877 => "0000000000000000",61878 => "0000000000000000",
61879 => "0000000000000000",61880 => "0000000000000000",
61881 => "0000000000000000",61882 => "0000000000000000",
61883 => "0000000000000000",61884 => "0000000000000000",
61885 => "0000000000000000",61886 => "0000000000000000",
61887 => "0000000000000000",61888 => "0000000000000000",
61889 => "0000000000000000",61890 => "0000000000000000",
61891 => "0000000000000000",61892 => "0000000000000000",
61893 => "0000000000000000",61894 => "0000000000000000",
61895 => "0000000000000000",61896 => "0000000000000000",
61897 => "0000000000000000",61898 => "0000000000000000",
61899 => "0000000000000000",61900 => "0000000000000000",
61901 => "0000000000000000",61902 => "0000000000000000",
61903 => "0000000000000000",61904 => "0000000000000000",
61905 => "0000000000000000",61906 => "0000000000000000",
61907 => "0000000000000000",61908 => "0000000000000000",
61909 => "0000000000000000",61910 => "0000000000000000",
61911 => "0000000000000000",61912 => "0000000000000000",
61913 => "0000000000000000",61914 => "0000000000000000",
61915 => "0000000000000000",61916 => "0000000000000000",
61917 => "0000000000000000",61918 => "0000000000000000",
61919 => "0000000000000000",61920 => "0000000000000000",
61921 => "0000000000000000",61922 => "0000000000000000",
61923 => "0000000000000000",61924 => "0000000000000000",
61925 => "0000000000000000",61926 => "0000000000000000",
61927 => "0000000000000000",61928 => "0000000000000000",
61929 => "0000000000000000",61930 => "0000000000000000",
61931 => "0000000000000000",61932 => "0000000000000000",
61933 => "0000000000000000",61934 => "0000000000000000",
61935 => "0000000000000000",61936 => "0000000000000000",
61937 => "0000000000000000",61938 => "0000000000000000",
61939 => "0000000000000000",61940 => "0000000000000000",
61941 => "0000000000000000",61942 => "0000000000000000",
61943 => "0000000000000000",61944 => "0000000000000000",
61945 => "0000000000000000",61946 => "0000000000000000",
61947 => "0000000000000000",61948 => "0000000000000000",
61949 => "0000000000000000",61950 => "0000000000000000",
61951 => "0000000000000000",61952 => "0000000000000000",
61953 => "0000000000000000",61954 => "0000000000000000",
61955 => "0000000000000000",61956 => "0000000000000000",
61957 => "0000000000000000",61958 => "0000000000000000",
61959 => "0000000000000000",61960 => "0000000000000000",
61961 => "0000000000000000",61962 => "0000000000000000",
61963 => "0000000000000000",61964 => "0000000000000000",
61965 => "0000000000000000",61966 => "0000000000000000",
61967 => "0000000000000000",61968 => "0000000000000000",
61969 => "0000000000000000",61970 => "0000000000000000",
61971 => "0000000000000000",61972 => "0000000000000000",
61973 => "0000000000000000",61974 => "0000000000000000",
61975 => "0000000000000000",61976 => "0000000000000000",
61977 => "0000000000000000",61978 => "0000000000000000",
61979 => "0000000000000000",61980 => "0000000000000000",
61981 => "0000000000000000",61982 => "0000000000000000",
61983 => "0000000000000000",61984 => "0000000000000000",
61985 => "0000000000000000",61986 => "0000000000000000",
61987 => "0000000000000000",61988 => "0000000000000000",
61989 => "0000000000000000",61990 => "0000000000000000",
61991 => "0000000000000000",61992 => "0000000000000000",
61993 => "0000000000000000",61994 => "0000000000000000",
61995 => "0000000000000000",61996 => "0000000000000000",
61997 => "0000000000000000",61998 => "0000000000000000",
61999 => "0000000000000000",62000 => "0000000000000000",
62001 => "0000000000000000",62002 => "0000000000000000",
62003 => "0000000000000000",62004 => "0000000000000000",
62005 => "0000000000000000",62006 => "0000000000000000",
62007 => "0000000000000000",62008 => "0000000000000000",
62009 => "0000000000000000",62010 => "0000000000000000",
62011 => "0000000000000000",62012 => "0000000000000000",
62013 => "0000000000000000",62014 => "0000000000000000",
62015 => "0000000000000000",62016 => "0000000000000000",
62017 => "0000000000000000",62018 => "0000000000000000",
62019 => "0000000000000000",62020 => "0000000000000000",
62021 => "0000000000000000",62022 => "0000000000000000",
62023 => "0000000000000000",62024 => "0000000000000000",
62025 => "0000000000000000",62026 => "0000000000000000",
62027 => "0000000000000000",62028 => "0000000000000000",
62029 => "0000000000000000",62030 => "0000000000000000",
62031 => "0000000000000000",62032 => "0000000000000000",
62033 => "0000000000000000",62034 => "0000000000000000",
62035 => "0000000000000000",62036 => "0000000000000000",
62037 => "0000000000000000",62038 => "0000000000000000",
62039 => "0000000000000000",62040 => "0000000000000000",
62041 => "0000000000000000",62042 => "0000000000000000",
62043 => "0000000000000000",62044 => "0000000000000000",
62045 => "0000000000000000",62046 => "0000000000000000",
62047 => "0000000000000000",62048 => "0000000000000000",
62049 => "0000000000000000",62050 => "0000000000000000",
62051 => "0000000000000000",62052 => "0000000000000000",
62053 => "0000000000000000",62054 => "0000000000000000",
62055 => "0000000000000000",62056 => "0000000000000000",
62057 => "0000000000000000",62058 => "0000000000000000",
62059 => "0000000000000000",62060 => "0000000000000000",
62061 => "0000000000000000",62062 => "0000000000000000",
62063 => "0000000000000000",62064 => "0000000000000000",
62065 => "0000000000000000",62066 => "0000000000000000",
62067 => "0000000000000000",62068 => "0000000000000000",
62069 => "0000000000000000",62070 => "0000000000000000",
62071 => "0000000000000000",62072 => "0000000000000000",
62073 => "0000000000000000",62074 => "0000000000000000",
62075 => "0000000000000000",62076 => "0000000000000000",
62077 => "0000000000000000",62078 => "0000000000000000",
62079 => "0000000000000000",62080 => "0000000000000000",
62081 => "0000000000000000",62082 => "0000000000000000",
62083 => "0000000000000000",62084 => "0000000000000000",
62085 => "0000000000000000",62086 => "0000000000000000",
62087 => "0000000000000000",62088 => "0000000000000000",
62089 => "0000000000000000",62090 => "0000000000000000",
62091 => "0000000000000000",62092 => "0000000000000000",
62093 => "0000000000000000",62094 => "0000000000000000",
62095 => "0000000000000000",62096 => "0000000000000000",
62097 => "0000000000000000",62098 => "0000000000000000",
62099 => "0000000000000000",62100 => "0000000000000000",
62101 => "0000000000000000",62102 => "0000000000000000",
62103 => "0000000000000000",62104 => "0000000000000000",
62105 => "0000000000000000",62106 => "0000000000000000",
62107 => "0000000000000000",62108 => "0000000000000000",
62109 => "0000000000000000",62110 => "0000000000000000",
62111 => "0000000000000000",62112 => "0000000000000000",
62113 => "0000000000000000",62114 => "0000000000000000",
62115 => "0000000000000000",62116 => "0000000000000000",
62117 => "0000000000000000",62118 => "0000000000000000",
62119 => "0000000000000000",62120 => "0000000000000000",
62121 => "0000000000000000",62122 => "0000000000000000",
62123 => "0000000000000000",62124 => "0000000000000000",
62125 => "0000000000000000",62126 => "0000000000000000",
62127 => "0000000000000000",62128 => "0000000000000000",
62129 => "0000000000000000",62130 => "0000000000000000",
62131 => "0000000000000000",62132 => "0000000000000000",
62133 => "0000000000000000",62134 => "0000000000000000",
62135 => "0000000000000000",62136 => "0000000000000000",
62137 => "0000000000000000",62138 => "0000000000000000",
62139 => "0000000000000000",62140 => "0000000000000000",
62141 => "0000000000000000",62142 => "0000000000000000",
62143 => "0000000000000000",62144 => "0000000000000000",
62145 => "0000000000000000",62146 => "0000000000000000",
62147 => "0000000000000000",62148 => "0000000000000000",
62149 => "0000000000000000",62150 => "0000000000000000",
62151 => "0000000000000000",62152 => "0000000000000000",
62153 => "0000000000000000",62154 => "0000000000000000",
62155 => "0000000000000000",62156 => "0000000000000000",
62157 => "0000000000000000",62158 => "0000000000000000",
62159 => "0000000000000000",62160 => "0000000000000000",
62161 => "0000000000000000",62162 => "0000000000000000",
62163 => "0000000000000000",62164 => "0000000000000000",
62165 => "0000000000000000",62166 => "0000000000000000",
62167 => "0000000000000000",62168 => "0000000000000000",
62169 => "0000000000000000",62170 => "0000000000000000",
62171 => "0000000000000000",62172 => "0000000000000000",
62173 => "0000000000000000",62174 => "0000000000000000",
62175 => "0000000000000000",62176 => "0000000000000000",
62177 => "0000000000000000",62178 => "0000000000000000",
62179 => "0000000000000000",62180 => "0000000000000000",
62181 => "0000000000000000",62182 => "0000000000000000",
62183 => "0000000000000000",62184 => "0000000000000000",
62185 => "0000000000000000",62186 => "0000000000000000",
62187 => "0000000000000000",62188 => "0000000000000000",
62189 => "0000000000000000",62190 => "0000000000000000",
62191 => "0000000000000000",62192 => "0000000000000000",
62193 => "0000000000000000",62194 => "0000000000000000",
62195 => "0000000000000000",62196 => "0000000000000000",
62197 => "0000000000000000",62198 => "0000000000000000",
62199 => "0000000000000000",62200 => "0000000000000000",
62201 => "0000000000000000",62202 => "0000000000000000",
62203 => "0000000000000000",62204 => "0000000000000000",
62205 => "0000000000000000",62206 => "0000000000000000",
62207 => "0000000000000000",62208 => "0000000000000000",
62209 => "0000000000000000",62210 => "0000000000000000",
62211 => "0000000000000000",62212 => "0000000000000000",
62213 => "0000000000000000",62214 => "0000000000000000",
62215 => "0000000000000000",62216 => "0000000000000000",
62217 => "0000000000000000",62218 => "0000000000000000",
62219 => "0000000000000000",62220 => "0000000000000000",
62221 => "0000000000000000",62222 => "0000000000000000",
62223 => "0000000000000000",62224 => "0000000000000000",
62225 => "0000000000000000",62226 => "0000000000000000",
62227 => "0000000000000000",62228 => "0000000000000000",
62229 => "0000000000000000",62230 => "0000000000000000",
62231 => "0000000000000000",62232 => "0000000000000000",
62233 => "0000000000000000",62234 => "0000000000000000",
62235 => "0000000000000000",62236 => "0000000000000000",
62237 => "0000000000000000",62238 => "0000000000000000",
62239 => "0000000000000000",62240 => "0000000000000000",
62241 => "0000000000000000",62242 => "0000000000000000",
62243 => "0000000000000000",62244 => "0000000000000000",
62245 => "0000000000000000",62246 => "0000000000000000",
62247 => "0000000000000000",62248 => "0000000000000000",
62249 => "0000000000000000",62250 => "0000000000000000",
62251 => "0000000000000000",62252 => "0000000000000000",
62253 => "0000000000000000",62254 => "0000000000000000",
62255 => "0000000000000000",62256 => "0000000000000000",
62257 => "0000000000000000",62258 => "0000000000000000",
62259 => "0000000000000000",62260 => "0000000000000000",
62261 => "0000000000000000",62262 => "0000000000000000",
62263 => "0000000000000000",62264 => "0000000000000000",
62265 => "0000000000000000",62266 => "0000000000000000",
62267 => "0000000000000000",62268 => "0000000000000000",
62269 => "0000000000000000",62270 => "0000000000000000",
62271 => "0000000000000000",62272 => "0000000000000000",
62273 => "0000000000000000",62274 => "0000000000000000",
62275 => "0000000000000000",62276 => "0000000000000000",
62277 => "0000000000000000",62278 => "0000000000000000",
62279 => "0000000000000000",62280 => "0000000000000000",
62281 => "0000000000000000",62282 => "0000000000000000",
62283 => "0000000000000000",62284 => "0000000000000000",
62285 => "0000000000000000",62286 => "0000000000000000",
62287 => "0000000000000000",62288 => "0000000000000000",
62289 => "0000000000000000",62290 => "0000000000000000",
62291 => "0000000000000000",62292 => "0000000000000000",
62293 => "0000000000000000",62294 => "0000000000000000",
62295 => "0000000000000000",62296 => "0000000000000000",
62297 => "0000000000000000",62298 => "0000000000000000",
62299 => "0000000000000000",62300 => "0000000000000000",
62301 => "0000000000000000",62302 => "0000000000000000",
62303 => "0000000000000000",62304 => "0000000000000000",
62305 => "0000000000000000",62306 => "0000000000000000",
62307 => "0000000000000000",62308 => "0000000000000000",
62309 => "0000000000000000",62310 => "0000000000000000",
62311 => "0000000000000000",62312 => "0000000000000000",
62313 => "0000000000000000",62314 => "0000000000000000",
62315 => "0000000000000000",62316 => "0000000000000000",
62317 => "0000000000000000",62318 => "0000000000000000",
62319 => "0000000000000000",62320 => "0000000000000000",
62321 => "0000000000000000",62322 => "0000000000000000",
62323 => "0000000000000000",62324 => "0000000000000000",
62325 => "0000000000000000",62326 => "0000000000000000",
62327 => "0000000000000000",62328 => "0000000000000000",
62329 => "0000000000000000",62330 => "0000000000000000",
62331 => "0000000000000000",62332 => "0000000000000000",
62333 => "0000000000000000",62334 => "0000000000000000",
62335 => "0000000000000000",62336 => "0000000000000000",
62337 => "0000000000000000",62338 => "0000000000000000",
62339 => "0000000000000000",62340 => "0000000000000000",
62341 => "0000000000000000",62342 => "0000000000000000",
62343 => "0000000000000000",62344 => "0000000000000000",
62345 => "0000000000000000",62346 => "0000000000000000",
62347 => "0000000000000000",62348 => "0000000000000000",
62349 => "0000000000000000",62350 => "0000000000000000",
62351 => "0000000000000000",62352 => "0000000000000000",
62353 => "0000000000000000",62354 => "0000000000000000",
62355 => "0000000000000000",62356 => "0000000000000000",
62357 => "0000000000000000",62358 => "0000000000000000",
62359 => "0000000000000000",62360 => "0000000000000000",
62361 => "0000000000000000",62362 => "0000000000000000",
62363 => "0000000000000000",62364 => "0000000000000000",
62365 => "0000000000000000",62366 => "0000000000000000",
62367 => "0000000000000000",62368 => "0000000000000000",
62369 => "0000000000000000",62370 => "0000000000000000",
62371 => "0000000000000000",62372 => "0000000000000000",
62373 => "0000000000000000",62374 => "0000000000000000",
62375 => "0000000000000000",62376 => "0000000000000000",
62377 => "0000000000000000",62378 => "0000000000000000",
62379 => "0000000000000000",62380 => "0000000000000000",
62381 => "0000000000000000",62382 => "0000000000000000",
62383 => "0000000000000000",62384 => "0000000000000000",
62385 => "0000000000000000",62386 => "0000000000000000",
62387 => "0000000000000000",62388 => "0000000000000000",
62389 => "0000000000000000",62390 => "0000000000000000",
62391 => "0000000000000000",62392 => "0000000000000000",
62393 => "0000000000000000",62394 => "0000000000000000",
62395 => "0000000000000000",62396 => "0000000000000000",
62397 => "0000000000000000",62398 => "0000000000000000",
62399 => "0000000000000000",62400 => "0000000000000000",
62401 => "0000000000000000",62402 => "0000000000000000",
62403 => "0000000000000000",62404 => "0000000000000000",
62405 => "0000000000000000",62406 => "0000000000000000",
62407 => "0000000000000000",62408 => "0000000000000000",
62409 => "0000000000000000",62410 => "0000000000000000",
62411 => "0000000000000000",62412 => "0000000000000000",
62413 => "0000000000000000",62414 => "0000000000000000",
62415 => "0000000000000000",62416 => "0000000000000000",
62417 => "0000000000000000",62418 => "0000000000000000",
62419 => "0000000000000000",62420 => "0000000000000000",
62421 => "0000000000000000",62422 => "0000000000000000",
62423 => "0000000000000000",62424 => "0000000000000000",
62425 => "0000000000000000",62426 => "0000000000000000",
62427 => "0000000000000000",62428 => "0000000000000000",
62429 => "0000000000000000",62430 => "0000000000000000",
62431 => "0000000000000000",62432 => "0000000000000000",
62433 => "0000000000000000",62434 => "0000000000000000",
62435 => "0000000000000000",62436 => "0000000000000000",
62437 => "0000000000000000",62438 => "0000000000000000",
62439 => "0000000000000000",62440 => "0000000000000000",
62441 => "0000000000000000",62442 => "0000000000000000",
62443 => "0000000000000000",62444 => "0000000000000000",
62445 => "0000000000000000",62446 => "0000000000000000",
62447 => "0000000000000000",62448 => "0000000000000000",
62449 => "0000000000000000",62450 => "0000000000000000",
62451 => "0000000000000000",62452 => "0000000000000000",
62453 => "0000000000000000",62454 => "0000000000000000",
62455 => "0000000000000000",62456 => "0000000000000000",
62457 => "0000000000000000",62458 => "0000000000000000",
62459 => "0000000000000000",62460 => "0000000000000000",
62461 => "0000000000000000",62462 => "0000000000000000",
62463 => "0000000000000000",62464 => "0000000000000000",
62465 => "0000000000000000",62466 => "0000000000000000",
62467 => "0000000000000000",62468 => "0000000000000000",
62469 => "0000000000000000",62470 => "0000000000000000",
62471 => "0000000000000000",62472 => "0000000000000000",
62473 => "0000000000000000",62474 => "0000000000000000",
62475 => "0000000000000000",62476 => "0000000000000000",
62477 => "0000000000000000",62478 => "0000000000000000",
62479 => "0000000000000000",62480 => "0000000000000000",
62481 => "0000000000000000",62482 => "0000000000000000",
62483 => "0000000000000000",62484 => "0000000000000000",
62485 => "0000000000000000",62486 => "0000000000000000",
62487 => "0000000000000000",62488 => "0000000000000000",
62489 => "0000000000000000",62490 => "0000000000000000",
62491 => "0000000000000000",62492 => "0000000000000000",
62493 => "0000000000000000",62494 => "0000000000000000",
62495 => "0000000000000000",62496 => "0000000000000000",
62497 => "0000000000000000",62498 => "0000000000000000",
62499 => "0000000000000000",62500 => "0000000000000000",
62501 => "0000000000000000",62502 => "0000000000000000",
62503 => "0000000000000000",62504 => "0000000000000000",
62505 => "0000000000000000",62506 => "0000000000000000",
62507 => "0000000000000000",62508 => "0000000000000000",
62509 => "0000000000000000",62510 => "0000000000000000",
62511 => "0000000000000000",62512 => "0000000000000000",
62513 => "0000000000000000",62514 => "0000000000000000",
62515 => "0000000000000000",62516 => "0000000000000000",
62517 => "0000000000000000",62518 => "0000000000000000",
62519 => "0000000000000000",62520 => "0000000000000000",
62521 => "0000000000000000",62522 => "0000000000000000",
62523 => "0000000000000000",62524 => "0000000000000000",
62525 => "0000000000000000",62526 => "0000000000000000",
62527 => "0000000000000000",62528 => "0000000000000000",
62529 => "0000000000000000",62530 => "0000000000000000",
62531 => "0000000000000000",62532 => "0000000000000000",
62533 => "0000000000000000",62534 => "0000000000000000",
62535 => "0000000000000000",62536 => "0000000000000000",
62537 => "0000000000000000",62538 => "0000000000000000",
62539 => "0000000000000000",62540 => "0000000000000000",
62541 => "0000000000000000",62542 => "0000000000000000",
62543 => "0000000000000000",62544 => "0000000000000000",
62545 => "0000000000000000",62546 => "0000000000000000",
62547 => "0000000000000000",62548 => "0000000000000000",
62549 => "0000000000000000",62550 => "0000000000000000",
62551 => "0000000000000000",62552 => "0000000000000000",
62553 => "0000000000000000",62554 => "0000000000000000",
62555 => "0000000000000000",62556 => "0000000000000000",
62557 => "0000000000000000",62558 => "0000000000000000",
62559 => "0000000000000000",62560 => "0000000000000000",
62561 => "0000000000000000",62562 => "0000000000000000",
62563 => "0000000000000000",62564 => "0000000000000000",
62565 => "0000000000000000",62566 => "0000000000000000",
62567 => "0000000000000000",62568 => "0000000000000000",
62569 => "0000000000000000",62570 => "0000000000000000",
62571 => "0000000000000000",62572 => "0000000000000000",
62573 => "0000000000000000",62574 => "0000000000000000",
62575 => "0000000000000000",62576 => "0000000000000000",
62577 => "0000000000000000",62578 => "0000000000000000",
62579 => "0000000000000000",62580 => "0000000000000000",
62581 => "0000000000000000",62582 => "0000000000000000",
62583 => "0000000000000000",62584 => "0000000000000000",
62585 => "0000000000000000",62586 => "0000000000000000",
62587 => "0000000000000000",62588 => "0000000000000000",
62589 => "0000000000000000",62590 => "0000000000000000",
62591 => "0000000000000000",62592 => "0000000000000000",
62593 => "0000000000000000",62594 => "0000000000000000",
62595 => "0000000000000000",62596 => "0000000000000000",
62597 => "0000000000000000",62598 => "0000000000000000",
62599 => "0000000000000000",62600 => "0000000000000000",
62601 => "0000000000000000",62602 => "0000000000000000",
62603 => "0000000000000000",62604 => "0000000000000000",
62605 => "0000000000000000",62606 => "0000000000000000",
62607 => "0000000000000000",62608 => "0000000000000000",
62609 => "0000000000000000",62610 => "0000000000000000",
62611 => "0000000000000000",62612 => "0000000000000000",
62613 => "0000000000000000",62614 => "0000000000000000",
62615 => "0000000000000000",62616 => "0000000000000000",
62617 => "0000000000000000",62618 => "0000000000000000",
62619 => "0000000000000000",62620 => "0000000000000000",
62621 => "0000000000000000",62622 => "0000000000000000",
62623 => "0000000000000000",62624 => "0000000000000000",
62625 => "0000000000000000",62626 => "0000000000000000",
62627 => "0000000000000000",62628 => "0000000000000000",
62629 => "0000000000000000",62630 => "0000000000000000",
62631 => "0000000000000000",62632 => "0000000000000000",
62633 => "0000000000000000",62634 => "0000000000000000",
62635 => "0000000000000000",62636 => "0000000000000000",
62637 => "0000000000000000",62638 => "0000000000000000",
62639 => "0000000000000000",62640 => "0000000000000000",
62641 => "0000000000000000",62642 => "0000000000000000",
62643 => "0000000000000000",62644 => "0000000000000000",
62645 => "0000000000000000",62646 => "0000000000000000",
62647 => "0000000000000000",62648 => "0000000000000000",
62649 => "0000000000000000",62650 => "0000000000000000",
62651 => "0000000000000000",62652 => "0000000000000000",
62653 => "0000000000000000",62654 => "0000000000000000",
62655 => "0000000000000000",62656 => "0000000000000000",
62657 => "0000000000000000",62658 => "0000000000000000",
62659 => "0000000000000000",62660 => "0000000000000000",
62661 => "0000000000000000",62662 => "0000000000000000",
62663 => "0000000000000000",62664 => "0000000000000000",
62665 => "0000000000000000",62666 => "0000000000000000",
62667 => "0000000000000000",62668 => "0000000000000000",
62669 => "0000000000000000",62670 => "0000000000000000",
62671 => "0000000000000000",62672 => "0000000000000000",
62673 => "0000000000000000",62674 => "0000000000000000",
62675 => "0000000000000000",62676 => "0000000000000000",
62677 => "0000000000000000",62678 => "0000000000000000",
62679 => "0000000000000000",62680 => "0000000000000000",
62681 => "0000000000000000",62682 => "0000000000000000",
62683 => "0000000000000000",62684 => "0000000000000000",
62685 => "0000000000000000",62686 => "0000000000000000",
62687 => "0000000000000000",62688 => "0000000000000000",
62689 => "0000000000000000",62690 => "0000000000000000",
62691 => "0000000000000000",62692 => "0000000000000000",
62693 => "0000000000000000",62694 => "0000000000000000",
62695 => "0000000000000000",62696 => "0000000000000000",
62697 => "0000000000000000",62698 => "0000000000000000",
62699 => "0000000000000000",62700 => "0000000000000000",
62701 => "0000000000000000",62702 => "0000000000000000",
62703 => "0000000000000000",62704 => "0000000000000000",
62705 => "0000000000000000",62706 => "0000000000000000",
62707 => "0000000000000000",62708 => "0000000000000000",
62709 => "0000000000000000",62710 => "0000000000000000",
62711 => "0000000000000000",62712 => "0000000000000000",
62713 => "0000000000000000",62714 => "0000000000000000",
62715 => "0000000000000000",62716 => "0000000000000000",
62717 => "0000000000000000",62718 => "0000000000000000",
62719 => "0000000000000000",62720 => "0000000000000000",
62721 => "0000000000000000",62722 => "0000000000000000",
62723 => "0000000000000000",62724 => "0000000000000000",
62725 => "0000000000000000",62726 => "0000000000000000",
62727 => "0000000000000000",62728 => "0000000000000000",
62729 => "0000000000000000",62730 => "0000000000000000",
62731 => "0000000000000000",62732 => "0000000000000000",
62733 => "0000000000000000",62734 => "0000000000000000",
62735 => "0000000000000000",62736 => "0000000000000000",
62737 => "0000000000000000",62738 => "0000000000000000",
62739 => "0000000000000000",62740 => "0000000000000000",
62741 => "0000000000000000",62742 => "0000000000000000",
62743 => "0000000000000000",62744 => "0000000000000000",
62745 => "0000000000000000",62746 => "0000000000000000",
62747 => "0000000000000000",62748 => "0000000000000000",
62749 => "0000000000000000",62750 => "0000000000000000",
62751 => "0000000000000000",62752 => "0000000000000000",
62753 => "0000000000000000",62754 => "0000000000000000",
62755 => "0000000000000000",62756 => "0000000000000000",
62757 => "0000000000000000",62758 => "0000000000000000",
62759 => "0000000000000000",62760 => "0000000000000000",
62761 => "0000000000000000",62762 => "0000000000000000",
62763 => "0000000000000000",62764 => "0000000000000000",
62765 => "0000000000000000",62766 => "0000000000000000",
62767 => "0000000000000000",62768 => "0000000000000000",
62769 => "0000000000000000",62770 => "0000000000000000",
62771 => "0000000000000000",62772 => "0000000000000000",
62773 => "0000000000000000",62774 => "0000000000000000",
62775 => "0000000000000000",62776 => "0000000000000000",
62777 => "0000000000000000",62778 => "0000000000000000",
62779 => "0000000000000000",62780 => "0000000000000000",
62781 => "0000000000000000",62782 => "0000000000000000",
62783 => "0000000000000000",62784 => "0000000000000000",
62785 => "0000000000000000",62786 => "0000000000000000",
62787 => "0000000000000000",62788 => "0000000000000000",
62789 => "0000000000000000",62790 => "0000000000000000",
62791 => "0000000000000000",62792 => "0000000000000000",
62793 => "0000000000000000",62794 => "0000000000000000",
62795 => "0000000000000000",62796 => "0000000000000000",
62797 => "0000000000000000",62798 => "0000000000000000",
62799 => "0000000000000000",62800 => "0000000000000000",
62801 => "0000000000000000",62802 => "0000000000000000",
62803 => "0000000000000000",62804 => "0000000000000000",
62805 => "0000000000000000",62806 => "0000000000000000",
62807 => "0000000000000000",62808 => "0000000000000000",
62809 => "0000000000000000",62810 => "0000000000000000",
62811 => "0000000000000000",62812 => "0000000000000000",
62813 => "0000000000000000",62814 => "0000000000000000",
62815 => "0000000000000000",62816 => "0000000000000000",
62817 => "0000000000000000",62818 => "0000000000000000",
62819 => "0000000000000000",62820 => "0000000000000000",
62821 => "0000000000000000",62822 => "0000000000000000",
62823 => "0000000000000000",62824 => "0000000000000000",
62825 => "0000000000000000",62826 => "0000000000000000",
62827 => "0000000000000000",62828 => "0000000000000000",
62829 => "0000000000000000",62830 => "0000000000000000",
62831 => "0000000000000000",62832 => "0000000000000000",
62833 => "0000000000000000",62834 => "0000000000000000",
62835 => "0000000000000000",62836 => "0000000000000000",
62837 => "0000000000000000",62838 => "0000000000000000",
62839 => "0000000000000000",62840 => "0000000000000000",
62841 => "0000000000000000",62842 => "0000000000000000",
62843 => "0000000000000000",62844 => "0000000000000000",
62845 => "0000000000000000",62846 => "0000000000000000",
62847 => "0000000000000000",62848 => "0000000000000000",
62849 => "0000000000000000",62850 => "0000000000000000",
62851 => "0000000000000000",62852 => "0000000000000000",
62853 => "0000000000000000",62854 => "0000000000000000",
62855 => "0000000000000000",62856 => "0000000000000000",
62857 => "0000000000000000",62858 => "0000000000000000",
62859 => "0000000000000000",62860 => "0000000000000000",
62861 => "0000000000000000",62862 => "0000000000000000",
62863 => "0000000000000000",62864 => "0000000000000000",
62865 => "0000000000000000",62866 => "0000000000000000",
62867 => "0000000000000000",62868 => "0000000000000000",
62869 => "0000000000000000",62870 => "0000000000000000",
62871 => "0000000000000000",62872 => "0000000000000000",
62873 => "0000000000000000",62874 => "0000000000000000",
62875 => "0000000000000000",62876 => "0000000000000000",
62877 => "0000000000000000",62878 => "0000000000000000",
62879 => "0000000000000000",62880 => "0000000000000000",
62881 => "0000000000000000",62882 => "0000000000000000",
62883 => "0000000000000000",62884 => "0000000000000000",
62885 => "0000000000000000",62886 => "0000000000000000",
62887 => "0000000000000000",62888 => "0000000000000000",
62889 => "0000000000000000",62890 => "0000000000000000",
62891 => "0000000000000000",62892 => "0000000000000000",
62893 => "0000000000000000",62894 => "0000000000000000",
62895 => "0000000000000000",62896 => "0000000000000000",
62897 => "0000000000000000",62898 => "0000000000000000",
62899 => "0000000000000000",62900 => "0000000000000000",
62901 => "0000000000000000",62902 => "0000000000000000",
62903 => "0000000000000000",62904 => "0000000000000000",
62905 => "0000000000000000",62906 => "0000000000000000",
62907 => "0000000000000000",62908 => "0000000000000000",
62909 => "0000000000000000",62910 => "0000000000000000",
62911 => "0000000000000000",62912 => "0000000000000000",
62913 => "0000000000000000",62914 => "0000000000000000",
62915 => "0000000000000000",62916 => "0000000000000000",
62917 => "0000000000000000",62918 => "0000000000000000",
62919 => "0000000000000000",62920 => "0000000000000000",
62921 => "0000000000000000",62922 => "0000000000000000",
62923 => "0000000000000000",62924 => "0000000000000000",
62925 => "0000000000000000",62926 => "0000000000000000",
62927 => "0000000000000000",62928 => "0000000000000000",
62929 => "0000000000000000",62930 => "0000000000000000",
62931 => "0000000000000000",62932 => "0000000000000000",
62933 => "0000000000000000",62934 => "0000000000000000",
62935 => "0000000000000000",62936 => "0000000000000000",
62937 => "0000000000000000",62938 => "0000000000000000",
62939 => "0000000000000000",62940 => "0000000000000000",
62941 => "0000000000000000",62942 => "0000000000000000",
62943 => "0000000000000000",62944 => "0000000000000000",
62945 => "0000000000000000",62946 => "0000000000000000",
62947 => "0000000000000000",62948 => "0000000000000000",
62949 => "0000000000000000",62950 => "0000000000000000",
62951 => "0000000000000000",62952 => "0000000000000000",
62953 => "0000000000000000",62954 => "0000000000000000",
62955 => "0000000000000000",62956 => "0000000000000000",
62957 => "0000000000000000",62958 => "0000000000000000",
62959 => "0000000000000000",62960 => "0000000000000000",
62961 => "0000000000000000",62962 => "0000000000000000",
62963 => "0000000000000000",62964 => "0000000000000000",
62965 => "0000000000000000",62966 => "0000000000000000",
62967 => "0000000000000000",62968 => "0000000000000000",
62969 => "0000000000000000",62970 => "0000000000000000",
62971 => "0000000000000000",62972 => "0000000000000000",
62973 => "0000000000000000",62974 => "0000000000000000",
62975 => "0000000000000000",62976 => "0000000000000000",
62977 => "0000000000000000",62978 => "0000000000000000",
62979 => "0000000000000000",62980 => "0000000000000000",
62981 => "0000000000000000",62982 => "0000000000000000",
62983 => "0000000000000000",62984 => "0000000000000000",
62985 => "0000000000000000",62986 => "0000000000000000",
62987 => "0000000000000000",62988 => "0000000000000000",
62989 => "0000000000000000",62990 => "0000000000000000",
62991 => "0000000000000000",62992 => "0000000000000000",
62993 => "0000000000000000",62994 => "0000000000000000",
62995 => "0000000000000000",62996 => "0000000000000000",
62997 => "0000000000000000",62998 => "0000000000000000",
62999 => "0000000000000000",63000 => "0000000000000000",
63001 => "0000000000000000",63002 => "0000000000000000",
63003 => "0000000000000000",63004 => "0000000000000000",
63005 => "0000000000000000",63006 => "0000000000000000",
63007 => "0000000000000000",63008 => "0000000000000000",
63009 => "0000000000000000",63010 => "0000000000000000",
63011 => "0000000000000000",63012 => "0000000000000000",
63013 => "0000000000000000",63014 => "0000000000000000",
63015 => "0000000000000000",63016 => "0000000000000000",
63017 => "0000000000000000",63018 => "0000000000000000",
63019 => "0000000000000000",63020 => "0000000000000000",
63021 => "0000000000000000",63022 => "0000000000000000",
63023 => "0000000000000000",63024 => "0000000000000000",
63025 => "0000000000000000",63026 => "0000000000000000",
63027 => "0000000000000000",63028 => "0000000000000000",
63029 => "0000000000000000",63030 => "0000000000000000",
63031 => "0000000000000000",63032 => "0000000000000000",
63033 => "0000000000000000",63034 => "0000000000000000",
63035 => "0000000000000000",63036 => "0000000000000000",
63037 => "0000000000000000",63038 => "0000000000000000",
63039 => "0000000000000000",63040 => "0000000000000000",
63041 => "0000000000000000",63042 => "0000000000000000",
63043 => "0000000000000000",63044 => "0000000000000000",
63045 => "0000000000000000",63046 => "0000000000000000",
63047 => "0000000000000000",63048 => "0000000000000000",
63049 => "0000000000000000",63050 => "0000000000000000",
63051 => "0000000000000000",63052 => "0000000000000000",
63053 => "0000000000000000",63054 => "0000000000000000",
63055 => "0000000000000000",63056 => "0000000000000000",
63057 => "0000000000000000",63058 => "0000000000000000",
63059 => "0000000000000000",63060 => "0000000000000000",
63061 => "0000000000000000",63062 => "0000000000000000",
63063 => "0000000000000000",63064 => "0000000000000000",
63065 => "0000000000000000",63066 => "0000000000000000",
63067 => "0000000000000000",63068 => "0000000000000000",
63069 => "0000000000000000",63070 => "0000000000000000",
63071 => "0000000000000000",63072 => "0000000000000000",
63073 => "0000000000000000",63074 => "0000000000000000",
63075 => "0000000000000000",63076 => "0000000000000000",
63077 => "0000000000000000",63078 => "0000000000000000",
63079 => "0000000000000000",63080 => "0000000000000000",
63081 => "0000000000000000",63082 => "0000000000000000",
63083 => "0000000000000000",63084 => "0000000000000000",
63085 => "0000000000000000",63086 => "0000000000000000",
63087 => "0000000000000000",63088 => "0000000000000000",
63089 => "0000000000000000",63090 => "0000000000000000",
63091 => "0000000000000000",63092 => "0000000000000000",
63093 => "0000000000000000",63094 => "0000000000000000",
63095 => "0000000000000000",63096 => "0000000000000000",
63097 => "0000000000000000",63098 => "0000000000000000",
63099 => "0000000000000000",63100 => "0000000000000000",
63101 => "0000000000000000",63102 => "0000000000000000",
63103 => "0000000000000000",63104 => "0000000000000000",
63105 => "0000000000000000",63106 => "0000000000000000",
63107 => "0000000000000000",63108 => "0000000000000000",
63109 => "0000000000000000",63110 => "0000000000000000",
63111 => "0000000000000000",63112 => "0000000000000000",
63113 => "0000000000000000",63114 => "0000000000000000",
63115 => "0000000000000000",63116 => "0000000000000000",
63117 => "0000000000000000",63118 => "0000000000000000",
63119 => "0000000000000000",63120 => "0000000000000000",
63121 => "0000000000000000",63122 => "0000000000000000",
63123 => "0000000000000000",63124 => "0000000000000000",
63125 => "0000000000000000",63126 => "0000000000000000",
63127 => "0000000000000000",63128 => "0000000000000000",
63129 => "0000000000000000",63130 => "0000000000000000",
63131 => "0000000000000000",63132 => "0000000000000000",
63133 => "0000000000000000",63134 => "0000000000000000",
63135 => "0000000000000000",63136 => "0000000000000000",
63137 => "0000000000000000",63138 => "0000000000000000",
63139 => "0000000000000000",63140 => "0000000000000000",
63141 => "0000000000000000",63142 => "0000000000000000",
63143 => "0000000000000000",63144 => "0000000000000000",
63145 => "0000000000000000",63146 => "0000000000000000",
63147 => "0000000000000000",63148 => "0000000000000000",
63149 => "0000000000000000",63150 => "0000000000000000",
63151 => "0000000000000000",63152 => "0000000000000000",
63153 => "0000000000000000",63154 => "0000000000000000",
63155 => "0000000000000000",63156 => "0000000000000000",
63157 => "0000000000000000",63158 => "0000000000000000",
63159 => "0000000000000000",63160 => "0000000000000000",
63161 => "0000000000000000",63162 => "0000000000000000",
63163 => "0000000000000000",63164 => "0000000000000000",
63165 => "0000000000000000",63166 => "0000000000000000",
63167 => "0000000000000000",63168 => "0000000000000000",
63169 => "0000000000000000",63170 => "0000000000000000",
63171 => "0000000000000000",63172 => "0000000000000000",
63173 => "0000000000000000",63174 => "0000000000000000",
63175 => "0000000000000000",63176 => "0000000000000000",
63177 => "0000000000000000",63178 => "0000000000000000",
63179 => "0000000000000000",63180 => "0000000000000000",
63181 => "0000000000000000",63182 => "0000000000000000",
63183 => "0000000000000000",63184 => "0000000000000000",
63185 => "0000000000000000",63186 => "0000000000000000",
63187 => "0000000000000000",63188 => "0000000000000000",
63189 => "0000000000000000",63190 => "0000000000000000",
63191 => "0000000000000000",63192 => "0000000000000000",
63193 => "0000000000000000",63194 => "0000000000000000",
63195 => "0000000000000000",63196 => "0000000000000000",
63197 => "0000000000000000",63198 => "0000000000000000",
63199 => "0000000000000000",63200 => "0000000000000000",
63201 => "0000000000000000",63202 => "0000000000000000",
63203 => "0000000000000000",63204 => "0000000000000000",
63205 => "0000000000000000",63206 => "0000000000000000",
63207 => "0000000000000000",63208 => "0000000000000000",
63209 => "0000000000000000",63210 => "0000000000000000",
63211 => "0000000000000000",63212 => "0000000000000000",
63213 => "0000000000000000",63214 => "0000000000000000",
63215 => "0000000000000000",63216 => "0000000000000000",
63217 => "0000000000000000",63218 => "0000000000000000",
63219 => "0000000000000000",63220 => "0000000000000000",
63221 => "0000000000000000",63222 => "0000000000000000",
63223 => "0000000000000000",63224 => "0000000000000000",
63225 => "0000000000000000",63226 => "0000000000000000",
63227 => "0000000000000000",63228 => "0000000000000000",
63229 => "0000000000000000",63230 => "0000000000000000",
63231 => "0000000000000000",63232 => "0000000000000000",
63233 => "0000000000000000",63234 => "0000000000000000",
63235 => "0000000000000000",63236 => "0000000000000000",
63237 => "0000000000000000",63238 => "0000000000000000",
63239 => "0000000000000000",63240 => "0000000000000000",
63241 => "0000000000000000",63242 => "0000000000000000",
63243 => "0000000000000000",63244 => "0000000000000000",
63245 => "0000000000000000",63246 => "0000000000000000",
63247 => "0000000000000000",63248 => "0000000000000000",
63249 => "0000000000000000",63250 => "0000000000000000",
63251 => "0000000000000000",63252 => "0000000000000000",
63253 => "0000000000000000",63254 => "0000000000000000",
63255 => "0000000000000000",63256 => "0000000000000000",
63257 => "0000000000000000",63258 => "0000000000000000",
63259 => "0000000000000000",63260 => "0000000000000000",
63261 => "0000000000000000",63262 => "0000000000000000",
63263 => "0000000000000000",63264 => "0000000000000000",
63265 => "0000000000000000",63266 => "0000000000000000",
63267 => "0000000000000000",63268 => "0000000000000000",
63269 => "0000000000000000",63270 => "0000000000000000",
63271 => "0000000000000000",63272 => "0000000000000000",
63273 => "0000000000000000",63274 => "0000000000000000",
63275 => "0000000000000000",63276 => "0000000000000000",
63277 => "0000000000000000",63278 => "0000000000000000",
63279 => "0000000000000000",63280 => "0000000000000000",
63281 => "0000000000000000",63282 => "0000000000000000",
63283 => "0000000000000000",63284 => "0000000000000000",
63285 => "0000000000000000",63286 => "0000000000000000",
63287 => "0000000000000000",63288 => "0000000000000000",
63289 => "0000000000000000",63290 => "0000000000000000",
63291 => "0000000000000000",63292 => "0000000000000000",
63293 => "0000000000000000",63294 => "0000000000000000",
63295 => "0000000000000000",63296 => "0000000000000000",
63297 => "0000000000000000",63298 => "0000000000000000",
63299 => "0000000000000000",63300 => "0000000000000000",
63301 => "0000000000000000",63302 => "0000000000000000",
63303 => "0000000000000000",63304 => "0000000000000000",
63305 => "0000000000000000",63306 => "0000000000000000",
63307 => "0000000000000000",63308 => "0000000000000000",
63309 => "0000000000000000",63310 => "0000000000000000",
63311 => "0000000000000000",63312 => "0000000000000000",
63313 => "0000000000000000",63314 => "0000000000000000",
63315 => "0000000000000000",63316 => "0000000000000000",
63317 => "0000000000000000",63318 => "0000000000000000",
63319 => "0000000000000000",63320 => "0000000000000000",
63321 => "0000000000000000",63322 => "0000000000000000",
63323 => "0000000000000000",63324 => "0000000000000000",
63325 => "0000000000000000",63326 => "0000000000000000",
63327 => "0000000000000000",63328 => "0000000000000000",
63329 => "0000000000000000",63330 => "0000000000000000",
63331 => "0000000000000000",63332 => "0000000000000000",
63333 => "0000000000000000",63334 => "0000000000000000",
63335 => "0000000000000000",63336 => "0000000000000000",
63337 => "0000000000000000",63338 => "0000000000000000",
63339 => "0000000000000000",63340 => "0000000000000000",
63341 => "0000000000000000",63342 => "0000000000000000",
63343 => "0000000000000000",63344 => "0000000000000000",
63345 => "0000000000000000",63346 => "0000000000000000",
63347 => "0000000000000000",63348 => "0000000000000000",
63349 => "0000000000000000",63350 => "0000000000000000",
63351 => "0000000000000000",63352 => "0000000000000000",
63353 => "0000000000000000",63354 => "0000000000000000",
63355 => "0000000000000000",63356 => "0000000000000000",
63357 => "0000000000000000",63358 => "0000000000000000",
63359 => "0000000000000000",63360 => "0000000000000000",
63361 => "0000000000000000",63362 => "0000000000000000",
63363 => "0000000000000000",63364 => "0000000000000000",
63365 => "0000000000000000",63366 => "0000000000000000",
63367 => "0000000000000000",63368 => "0000000000000000",
63369 => "0000000000000000",63370 => "0000000000000000",
63371 => "0000000000000000",63372 => "0000000000000000",
63373 => "0000000000000000",63374 => "0000000000000000",
63375 => "0000000000000000",63376 => "0000000000000000",
63377 => "0000000000000000",63378 => "0000000000000000",
63379 => "0000000000000000",63380 => "0000000000000000",
63381 => "0000000000000000",63382 => "0000000000000000",
63383 => "0000000000000000",63384 => "0000000000000000",
63385 => "0000000000000000",63386 => "0000000000000000",
63387 => "0000000000000000",63388 => "0000000000000000",
63389 => "0000000000000000",63390 => "0000000000000000",
63391 => "0000000000000000",63392 => "0000000000000000",
63393 => "0000000000000000",63394 => "0000000000000000",
63395 => "0000000000000000",63396 => "0000000000000000",
63397 => "0000000000000000",63398 => "0000000000000000",
63399 => "0000000000000000",63400 => "0000000000000000",
63401 => "0000000000000000",63402 => "0000000000000000",
63403 => "0000000000000000",63404 => "0000000000000000",
63405 => "0000000000000000",63406 => "0000000000000000",
63407 => "0000000000000000",63408 => "0000000000000000",
63409 => "0000000000000000",63410 => "0000000000000000",
63411 => "0000000000000000",63412 => "0000000000000000",
63413 => "0000000000000000",63414 => "0000000000000000",
63415 => "0000000000000000",63416 => "0000000000000000",
63417 => "0000000000000000",63418 => "0000000000000000",
63419 => "0000000000000000",63420 => "0000000000000000",
63421 => "0000000000000000",63422 => "0000000000000000",
63423 => "0000000000000000",63424 => "0000000000000000",
63425 => "0000000000000000",63426 => "0000000000000000",
63427 => "0000000000000000",63428 => "0000000000000000",
63429 => "0000000000000000",63430 => "0000000000000000",
63431 => "0000000000000000",63432 => "0000000000000000",
63433 => "0000000000000000",63434 => "0000000000000000",
63435 => "0000000000000000",63436 => "0000000000000000",
63437 => "0000000000000000",63438 => "0000000000000000",
63439 => "0000000000000000",63440 => "0000000000000000",
63441 => "0000000000000000",63442 => "0000000000000000",
63443 => "0000000000000000",63444 => "0000000000000000",
63445 => "0000000000000000",63446 => "0000000000000000",
63447 => "0000000000000000",63448 => "0000000000000000",
63449 => "0000000000000000",63450 => "0000000000000000",
63451 => "0000000000000000",63452 => "0000000000000000",
63453 => "0000000000000000",63454 => "0000000000000000",
63455 => "0000000000000000",63456 => "0000000000000000",
63457 => "0000000000000000",63458 => "0000000000000000",
63459 => "0000000000000000",63460 => "0000000000000000",
63461 => "0000000000000000",63462 => "0000000000000000",
63463 => "0000000000000000",63464 => "0000000000000000",
63465 => "0000000000000000",63466 => "0000000000000000",
63467 => "0000000000000000",63468 => "0000000000000000",
63469 => "0000000000000000",63470 => "0000000000000000",
63471 => "0000000000000000",63472 => "0000000000000000",
63473 => "0000000000000000",63474 => "0000000000000000",
63475 => "0000000000000000",63476 => "0000000000000000",
63477 => "0000000000000000",63478 => "0000000000000000",
63479 => "0000000000000000",63480 => "0000000000000000",
63481 => "0000000000000000",63482 => "0000000000000000",
63483 => "0000000000000000",63484 => "0000000000000000",
63485 => "0000000000000000",63486 => "0000000000000000",
63487 => "0000000000000000",63488 => "0000000000000000",
63489 => "0000000000000000",63490 => "0000000000000000",
63491 => "0000000000000000",63492 => "0000000000000000",
63493 => "0000000000000000",63494 => "0000000000000000",
63495 => "0000000000000000",63496 => "0000000000000000",
63497 => "0000000000000000",63498 => "0000000000000000",
63499 => "0000000000000000",63500 => "0000000000000000",
63501 => "0000000000000000",63502 => "0000000000000000",
63503 => "0000000000000000",63504 => "0000000000000000",
63505 => "0000000000000000",63506 => "0000000000000000",
63507 => "0000000000000000",63508 => "0000000000000000",
63509 => "0000000000000000",63510 => "0000000000000000",
63511 => "0000000000000000",63512 => "0000000000000000",
63513 => "0000000000000000",63514 => "0000000000000000",
63515 => "0000000000000000",63516 => "0000000000000000",
63517 => "0000000000000000",63518 => "0000000000000000",
63519 => "0000000000000000",63520 => "0000000000000000",
63521 => "0000000000000000",63522 => "0000000000000000",
63523 => "0000000000000000",63524 => "0000000000000000",
63525 => "0000000000000000",63526 => "0000000000000000",
63527 => "0000000000000000",63528 => "0000000000000000",
63529 => "0000000000000000",63530 => "0000000000000000",
63531 => "0000000000000000",63532 => "0000000000000000",
63533 => "0000000000000000",63534 => "0000000000000000",
63535 => "0000000000000000",63536 => "0000000000000000",
63537 => "0000000000000000",63538 => "0000000000000000",
63539 => "0000000000000000",63540 => "0000000000000000",
63541 => "0000000000000000",63542 => "0000000000000000",
63543 => "0000000000000000",63544 => "0000000000000000",
63545 => "0000000000000000",63546 => "0000000000000000",
63547 => "0000000000000000",63548 => "0000000000000000",
63549 => "0000000000000000",63550 => "0000000000000000",
63551 => "0000000000000000",63552 => "0000000000000000",
63553 => "0000000000000000",63554 => "0000000000000000",
63555 => "0000000000000000",63556 => "0000000000000000",
63557 => "0000000000000000",63558 => "0000000000000000",
63559 => "0000000000000000",63560 => "0000000000000000",
63561 => "0000000000000000",63562 => "0000000000000000",
63563 => "0000000000000000",63564 => "0000000000000000",
63565 => "0000000000000000",63566 => "0000000000000000",
63567 => "0000000000000000",63568 => "0000000000000000",
63569 => "0000000000000000",63570 => "0000000000000000",
63571 => "0000000000000000",63572 => "0000000000000000",
63573 => "0000000000000000",63574 => "0000000000000000",
63575 => "0000000000000000",63576 => "0000000000000000",
63577 => "0000000000000000",63578 => "0000000000000000",
63579 => "0000000000000000",63580 => "0000000000000000",
63581 => "0000000000000000",63582 => "0000000000000000",
63583 => "0000000000000000",63584 => "0000000000000000",
63585 => "0000000000000000",63586 => "0000000000000000",
63587 => "0000000000000000",63588 => "0000000000000000",
63589 => "0000000000000000",63590 => "0000000000000000",
63591 => "0000000000000000",63592 => "0000000000000000",
63593 => "0000000000000000",63594 => "0000000000000000",
63595 => "0000000000000000",63596 => "0000000000000000",
63597 => "0000000000000000",63598 => "0000000000000000",
63599 => "0000000000000000",63600 => "0000000000000000",
63601 => "0000000000000000",63602 => "0000000000000000",
63603 => "0000000000000000",63604 => "0000000000000000",
63605 => "0000000000000000",63606 => "0000000000000000",
63607 => "0000000000000000",63608 => "0000000000000000",
63609 => "0000000000000000",63610 => "0000000000000000",
63611 => "0000000000000000",63612 => "0000000000000000",
63613 => "0000000000000000",63614 => "0000000000000000",
63615 => "0000000000000000",63616 => "0000000000000000",
63617 => "0000000000000000",63618 => "0000000000000000",
63619 => "0000000000000000",63620 => "0000000000000000",
63621 => "0000000000000000",63622 => "0000000000000000",
63623 => "0000000000000000",63624 => "0000000000000000",
63625 => "0000000000000000",63626 => "0000000000000000",
63627 => "0000000000000000",63628 => "0000000000000000",
63629 => "0000000000000000",63630 => "0000000000000000",
63631 => "0000000000000000",63632 => "0000000000000000",
63633 => "0000000000000000",63634 => "0000000000000000",
63635 => "0000000000000000",63636 => "0000000000000000",
63637 => "0000000000000000",63638 => "0000000000000000",
63639 => "0000000000000000",63640 => "0000000000000000",
63641 => "0000000000000000",63642 => "0000000000000000",
63643 => "0000000000000000",63644 => "0000000000000000",
63645 => "0000000000000000",63646 => "0000000000000000",
63647 => "0000000000000000",63648 => "0000000000000000",
63649 => "0000000000000000",63650 => "0000000000000000",
63651 => "0000000000000000",63652 => "0000000000000000",
63653 => "0000000000000000",63654 => "0000000000000000",
63655 => "0000000000000000",63656 => "0000000000000000",
63657 => "0000000000000000",63658 => "0000000000000000",
63659 => "0000000000000000",63660 => "0000000000000000",
63661 => "0000000000000000",63662 => "0000000000000000",
63663 => "0000000000000000",63664 => "0000000000000000",
63665 => "0000000000000000",63666 => "0000000000000000",
63667 => "0000000000000000",63668 => "0000000000000000",
63669 => "0000000000000000",63670 => "0000000000000000",
63671 => "0000000000000000",63672 => "0000000000000000",
63673 => "0000000000000000",63674 => "0000000000000000",
63675 => "0000000000000000",63676 => "0000000000000000",
63677 => "0000000000000000",63678 => "0000000000000000",
63679 => "0000000000000000",63680 => "0000000000000000",
63681 => "0000000000000000",63682 => "0000000000000000",
63683 => "0000000000000000",63684 => "0000000000000000",
63685 => "0000000000000000",63686 => "0000000000000000",
63687 => "0000000000000000",63688 => "0000000000000000",
63689 => "0000000000000000",63690 => "0000000000000000",
63691 => "0000000000000000",63692 => "0000000000000000",
63693 => "0000000000000000",63694 => "0000000000000000",
63695 => "0000000000000000",63696 => "0000000000000000",
63697 => "0000000000000000",63698 => "0000000000000000",
63699 => "0000000000000000",63700 => "0000000000000000",
63701 => "0000000000000000",63702 => "0000000000000000",
63703 => "0000000000000000",63704 => "0000000000000000",
63705 => "0000000000000000",63706 => "0000000000000000",
63707 => "0000000000000000",63708 => "0000000000000000",
63709 => "0000000000000000",63710 => "0000000000000000",
63711 => "0000000000000000",63712 => "0000000000000000",
63713 => "0000000000000000",63714 => "0000000000000000",
63715 => "0000000000000000",63716 => "0000000000000000",
63717 => "0000000000000000",63718 => "0000000000000000",
63719 => "0000000000000000",63720 => "0000000000000000",
63721 => "0000000000000000",63722 => "0000000000000000",
63723 => "0000000000000000",63724 => "0000000000000000",
63725 => "0000000000000000",63726 => "0000000000000000",
63727 => "0000000000000000",63728 => "0000000000000000",
63729 => "0000000000000000",63730 => "0000000000000000",
63731 => "0000000000000000",63732 => "0000000000000000",
63733 => "0000000000000000",63734 => "0000000000000000",
63735 => "0000000000000000",63736 => "0000000000000000",
63737 => "0000000000000000",63738 => "0000000000000000",
63739 => "0000000000000000",63740 => "0000000000000000",
63741 => "0000000000000000",63742 => "0000000000000000",
63743 => "0000000000000000",63744 => "0000000000000000",
63745 => "0000000000000000",63746 => "0000000000000000",
63747 => "0000000000000000",63748 => "0000000000000000",
63749 => "0000000000000000",63750 => "0000000000000000",
63751 => "0000000000000000",63752 => "0000000000000000",
63753 => "0000000000000000",63754 => "0000000000000000",
63755 => "0000000000000000",63756 => "0000000000000000",
63757 => "0000000000000000",63758 => "0000000000000000",
63759 => "0000000000000000",63760 => "0000000000000000",
63761 => "0000000000000000",63762 => "0000000000000000",
63763 => "0000000000000000",63764 => "0000000000000000",
63765 => "0000000000000000",63766 => "0000000000000000",
63767 => "0000000000000000",63768 => "0000000000000000",
63769 => "0000000000000000",63770 => "0000000000000000",
63771 => "0000000000000000",63772 => "0000000000000000",
63773 => "0000000000000000",63774 => "0000000000000000",
63775 => "0000000000000000",63776 => "0000000000000000",
63777 => "0000000000000000",63778 => "0000000000000000",
63779 => "0000000000000000",63780 => "0000000000000000",
63781 => "0000000000000000",63782 => "0000000000000000",
63783 => "0000000000000000",63784 => "0000000000000000",
63785 => "0000000000000000",63786 => "0000000000000000",
63787 => "0000000000000000",63788 => "0000000000000000",
63789 => "0000000000000000",63790 => "0000000000000000",
63791 => "0000000000000000",63792 => "0000000000000000",
63793 => "0000000000000000",63794 => "0000000000000000",
63795 => "0000000000000000",63796 => "0000000000000000",
63797 => "0000000000000000",63798 => "0000000000000000",
63799 => "0000000000000000",63800 => "0000000000000000",
63801 => "0000000000000000",63802 => "0000000000000000",
63803 => "0000000000000000",63804 => "0000000000000000",
63805 => "0000000000000000",63806 => "0000000000000000",
63807 => "0000000000000000",63808 => "0000000000000000",
63809 => "0000000000000000",63810 => "0000000000000000",
63811 => "0000000000000000",63812 => "0000000000000000",
63813 => "0000000000000000",63814 => "0000000000000000",
63815 => "0000000000000000",63816 => "0000000000000000",
63817 => "0000000000000000",63818 => "0000000000000000",
63819 => "0000000000000000",63820 => "0000000000000000",
63821 => "0000000000000000",63822 => "0000000000000000",
63823 => "0000000000000000",63824 => "0000000000000000",
63825 => "0000000000000000",63826 => "0000000000000000",
63827 => "0000000000000000",63828 => "0000000000000000",
63829 => "0000000000000000",63830 => "0000000000000000",
63831 => "0000000000000000",63832 => "0000000000000000",
63833 => "0000000000000000",63834 => "0000000000000000",
63835 => "0000000000000000",63836 => "0000000000000000",
63837 => "0000000000000000",63838 => "0000000000000000",
63839 => "0000000000000000",63840 => "0000000000000000",
63841 => "0000000000000000",63842 => "0000000000000000",
63843 => "0000000000000000",63844 => "0000000000000000",
63845 => "0000000000000000",63846 => "0000000000000000",
63847 => "0000000000000000",63848 => "0000000000000000",
63849 => "0000000000000000",63850 => "0000000000000000",
63851 => "0000000000000000",63852 => "0000000000000000",
63853 => "0000000000000000",63854 => "0000000000000000",
63855 => "0000000000000000",63856 => "0000000000000000",
63857 => "0000000000000000",63858 => "0000000000000000",
63859 => "0000000000000000",63860 => "0000000000000000",
63861 => "0000000000000000",63862 => "0000000000000000",
63863 => "0000000000000000",63864 => "0000000000000000",
63865 => "0000000000000000",63866 => "0000000000000000",
63867 => "0000000000000000",63868 => "0000000000000000",
63869 => "0000000000000000",63870 => "0000000000000000",
63871 => "0000000000000000",63872 => "0000000000000000",
63873 => "0000000000000000",63874 => "0000000000000000",
63875 => "0000000000000000",63876 => "0000000000000000",
63877 => "0000000000000000",63878 => "0000000000000000",
63879 => "0000000000000000",63880 => "0000000000000000",
63881 => "0000000000000000",63882 => "0000000000000000",
63883 => "0000000000000000",63884 => "0000000000000000",
63885 => "0000000000000000",63886 => "0000000000000000",
63887 => "0000000000000000",63888 => "0000000000000000",
63889 => "0000000000000000",63890 => "0000000000000000",
63891 => "0000000000000000",63892 => "0000000000000000",
63893 => "0000000000000000",63894 => "0000000000000000",
63895 => "0000000000000000",63896 => "0000000000000000",
63897 => "0000000000000000",63898 => "0000000000000000",
63899 => "0000000000000000",63900 => "0000000000000000",
63901 => "0000000000000000",63902 => "0000000000000000",
63903 => "0000000000000000",63904 => "0000000000000000",
63905 => "0000000000000000",63906 => "0000000000000000",
63907 => "0000000000000000",63908 => "0000000000000000",
63909 => "0000000000000000",63910 => "0000000000000000",
63911 => "0000000000000000",63912 => "0000000000000000",
63913 => "0000000000000000",63914 => "0000000000000000",
63915 => "0000000000000000",63916 => "0000000000000000",
63917 => "0000000000000000",63918 => "0000000000000000",
63919 => "0000000000000000",63920 => "0000000000000000",
63921 => "0000000000000000",63922 => "0000000000000000",
63923 => "0000000000000000",63924 => "0000000000000000",
63925 => "0000000000000000",63926 => "0000000000000000",
63927 => "0000000000000000",63928 => "0000000000000000",
63929 => "0000000000000000",63930 => "0000000000000000",
63931 => "0000000000000000",63932 => "0000000000000000",
63933 => "0000000000000000",63934 => "0000000000000000",
63935 => "0000000000000000",63936 => "0000000000000000",
63937 => "0000000000000000",63938 => "0000000000000000",
63939 => "0000000000000000",63940 => "0000000000000000",
63941 => "0000000000000000",63942 => "0000000000000000",
63943 => "0000000000000000",63944 => "0000000000000000",
63945 => "0000000000000000",63946 => "0000000000000000",
63947 => "0000000000000000",63948 => "0000000000000000",
63949 => "0000000000000000",63950 => "0000000000000000",
63951 => "0000000000000000",63952 => "0000000000000000",
63953 => "0000000000000000",63954 => "0000000000000000",
63955 => "0000000000000000",63956 => "0000000000000000",
63957 => "0000000000000000",63958 => "0000000000000000",
63959 => "0000000000000000",63960 => "0000000000000000",
63961 => "0000000000000000",63962 => "0000000000000000",
63963 => "0000000000000000",63964 => "0000000000000000",
63965 => "0000000000000000",63966 => "0000000000000000",
63967 => "0000000000000000",63968 => "0000000000000000",
63969 => "0000000000000000",63970 => "0000000000000000",
63971 => "0000000000000000",63972 => "0000000000000000",
63973 => "0000000000000000",63974 => "0000000000000000",
63975 => "0000000000000000",63976 => "0000000000000000",
63977 => "0000000000000000",63978 => "0000000000000000",
63979 => "0000000000000000",63980 => "0000000000000000",
63981 => "0000000000000000",63982 => "0000000000000000",
63983 => "0000000000000000",63984 => "0000000000000000",
63985 => "0000000000000000",63986 => "0000000000000000",
63987 => "0000000000000000",63988 => "0000000000000000",
63989 => "0000000000000000",63990 => "0000000000000000",
63991 => "0000000000000000",63992 => "0000000000000000",
63993 => "0000000000000000",63994 => "0000000000000000",
63995 => "0000000000000000",63996 => "0000000000000000",
63997 => "0000000000000000",63998 => "0000000000000000",
63999 => "0000000000000000",64000 => "0000000000000000",
64001 => "0000000000000000",64002 => "0000000000000000",
64003 => "0000000000000000",64004 => "0000000000000000",
64005 => "0000000000000000",64006 => "0000000000000000",
64007 => "0000000000000000",64008 => "0000000000000000",
64009 => "0000000000000000",64010 => "0000000000000000",
64011 => "0000000000000000",64012 => "0000000000000000",
64013 => "0000000000000000",64014 => "0000000000000000",
64015 => "0000000000000000",64016 => "0000000000000000",
64017 => "0000000000000000",64018 => "0000000000000000",
64019 => "0000000000000000",64020 => "0000000000000000",
64021 => "0000000000000000",64022 => "0000000000000000",
64023 => "0000000000000000",64024 => "0000000000000000",
64025 => "0000000000000000",64026 => "0000000000000000",
64027 => "0000000000000000",64028 => "0000000000000000",
64029 => "0000000000000000",64030 => "0000000000000000",
64031 => "0000000000000000",64032 => "0000000000000000",
64033 => "0000000000000000",64034 => "0000000000000000",
64035 => "0000000000000000",64036 => "0000000000000000",
64037 => "0000000000000000",64038 => "0000000000000000",
64039 => "0000000000000000",64040 => "0000000000000000",
64041 => "0000000000000000",64042 => "0000000000000000",
64043 => "0000000000000000",64044 => "0000000000000000",
64045 => "0000000000000000",64046 => "0000000000000000",
64047 => "0000000000000000",64048 => "0000000000000000",
64049 => "0000000000000000",64050 => "0000000000000000",
64051 => "0000000000000000",64052 => "0000000000000000",
64053 => "0000000000000000",64054 => "0000000000000000",
64055 => "0000000000000000",64056 => "0000000000000000",
64057 => "0000000000000000",64058 => "0000000000000000",
64059 => "0000000000000000",64060 => "0000000000000000",
64061 => "0000000000000000",64062 => "0000000000000000",
64063 => "0000000000000000",64064 => "0000000000000000",
64065 => "0000000000000000",64066 => "0000000000000000",
64067 => "0000000000000000",64068 => "0000000000000000",
64069 => "0000000000000000",64070 => "0000000000000000",
64071 => "0000000000000000",64072 => "0000000000000000",
64073 => "0000000000000000",64074 => "0000000000000000",
64075 => "0000000000000000",64076 => "0000000000000000",
64077 => "0000000000000000",64078 => "0000000000000000",
64079 => "0000000000000000",64080 => "0000000000000000",
64081 => "0000000000000000",64082 => "0000000000000000",
64083 => "0000000000000000",64084 => "0000000000000000",
64085 => "0000000000000000",64086 => "0000000000000000",
64087 => "0000000000000000",64088 => "0000000000000000",
64089 => "0000000000000000",64090 => "0000000000000000",
64091 => "0000000000000000",64092 => "0000000000000000",
64093 => "0000000000000000",64094 => "0000000000000000",
64095 => "0000000000000000",64096 => "0000000000000000",
64097 => "0000000000000000",64098 => "0000000000000000",
64099 => "0000000000000000",64100 => "0000000000000000",
64101 => "0000000000000000",64102 => "0000000000000000",
64103 => "0000000000000000",64104 => "0000000000000000",
64105 => "0000000000000000",64106 => "0000000000000000",
64107 => "0000000000000000",64108 => "0000000000000000",
64109 => "0000000000000000",64110 => "0000000000000000",
64111 => "0000000000000000",64112 => "0000000000000000",
64113 => "0000000000000000",64114 => "0000000000000000",
64115 => "0000000000000000",64116 => "0000000000000000",
64117 => "0000000000000000",64118 => "0000000000000000",
64119 => "0000000000000000",64120 => "0000000000000000",
64121 => "0000000000000000",64122 => "0000000000000000",
64123 => "0000000000000000",64124 => "0000000000000000",
64125 => "0000000000000000",64126 => "0000000000000000",
64127 => "0000000000000000",64128 => "0000000000000000",
64129 => "0000000000000000",64130 => "0000000000000000",
64131 => "0000000000000000",64132 => "0000000000000000",
64133 => "0000000000000000",64134 => "0000000000000000",
64135 => "0000000000000000",64136 => "0000000000000000",
64137 => "0000000000000000",64138 => "0000000000000000",
64139 => "0000000000000000",64140 => "0000000000000000",
64141 => "0000000000000000",64142 => "0000000000000000",
64143 => "0000000000000000",64144 => "0000000000000000",
64145 => "0000000000000000",64146 => "0000000000000000",
64147 => "0000000000000000",64148 => "0000000000000000",
64149 => "0000000000000000",64150 => "0000000000000000",
64151 => "0000000000000000",64152 => "0000000000000000",
64153 => "0000000000000000",64154 => "0000000000000000",
64155 => "0000000000000000",64156 => "0000000000000000",
64157 => "0000000000000000",64158 => "0000000000000000",
64159 => "0000000000000000",64160 => "0000000000000000",
64161 => "0000000000000000",64162 => "0000000000000000",
64163 => "0000000000000000",64164 => "0000000000000000",
64165 => "0000000000000000",64166 => "0000000000000000",
64167 => "0000000000000000",64168 => "0000000000000000",
64169 => "0000000000000000",64170 => "0000000000000000",
64171 => "0000000000000000",64172 => "0000000000000000",
64173 => "0000000000000000",64174 => "0000000000000000",
64175 => "0000000000000000",64176 => "0000000000000000",
64177 => "0000000000000000",64178 => "0000000000000000",
64179 => "0000000000000000",64180 => "0000000000000000",
64181 => "0000000000000000",64182 => "0000000000000000",
64183 => "0000000000000000",64184 => "0000000000000000",
64185 => "0000000000000000",64186 => "0000000000000000",
64187 => "0000000000000000",64188 => "0000000000000000",
64189 => "0000000000000000",64190 => "0000000000000000",
64191 => "0000000000000000",64192 => "0000000000000000",
64193 => "0000000000000000",64194 => "0000000000000000",
64195 => "0000000000000000",64196 => "0000000000000000",
64197 => "0000000000000000",64198 => "0000000000000000",
64199 => "0000000000000000",64200 => "0000000000000000",
64201 => "0000000000000000",64202 => "0000000000000000",
64203 => "0000000000000000",64204 => "0000000000000000",
64205 => "0000000000000000",64206 => "0000000000000000",
64207 => "0000000000000000",64208 => "0000000000000000",
64209 => "0000000000000000",64210 => "0000000000000000",
64211 => "0000000000000000",64212 => "0000000000000000",
64213 => "0000000000000000",64214 => "0000000000000000",
64215 => "0000000000000000",64216 => "0000000000000000",
64217 => "0000000000000000",64218 => "0000000000000000",
64219 => "0000000000000000",64220 => "0000000000000000",
64221 => "0000000000000000",64222 => "0000000000000000",
64223 => "0000000000000000",64224 => "0000000000000000",
64225 => "0000000000000000",64226 => "0000000000000000",
64227 => "0000000000000000",64228 => "0000000000000000",
64229 => "0000000000000000",64230 => "0000000000000000",
64231 => "0000000000000000",64232 => "0000000000000000",
64233 => "0000000000000000",64234 => "0000000000000000",
64235 => "0000000000000000",64236 => "0000000000000000",
64237 => "0000000000000000",64238 => "0000000000000000",
64239 => "0000000000000000",64240 => "0000000000000000",
64241 => "0000000000000000",64242 => "0000000000000000",
64243 => "0000000000000000",64244 => "0000000000000000",
64245 => "0000000000000000",64246 => "0000000000000000",
64247 => "0000000000000000",64248 => "0000000000000000",
64249 => "0000000000000000",64250 => "0000000000000000",
64251 => "0000000000000000",64252 => "0000000000000000",
64253 => "0000000000000000",64254 => "0000000000000000",
64255 => "0000000000000000",64256 => "0000000000000000",
64257 => "0000000000000000",64258 => "0000000000000000",
64259 => "0000000000000000",64260 => "0000000000000000",
64261 => "0000000000000000",64262 => "0000000000000000",
64263 => "0000000000000000",64264 => "0000000000000000",
64265 => "0000000000000000",64266 => "0000000000000000",
64267 => "0000000000000000",64268 => "0000000000000000",
64269 => "0000000000000000",64270 => "0000000000000000",
64271 => "0000000000000000",64272 => "0000000000000000",
64273 => "0000000000000000",64274 => "0000000000000000",
64275 => "0000000000000000",64276 => "0000000000000000",
64277 => "0000000000000000",64278 => "0000000000000000",
64279 => "0000000000000000",64280 => "0000000000000000",
64281 => "0000000000000000",64282 => "0000000000000000",
64283 => "0000000000000000",64284 => "0000000000000000",
64285 => "0000000000000000",64286 => "0000000000000000",
64287 => "0000000000000000",64288 => "0000000000000000",
64289 => "0000000000000000",64290 => "0000000000000000",
64291 => "0000000000000000",64292 => "0000000000000000",
64293 => "0000000000000000",64294 => "0000000000000000",
64295 => "0000000000000000",64296 => "0000000000000000",
64297 => "0000000000000000",64298 => "0000000000000000",
64299 => "0000000000000000",64300 => "0000000000000000",
64301 => "0000000000000000",64302 => "0000000000000000",
64303 => "0000000000000000",64304 => "0000000000000000",
64305 => "0000000000000000",64306 => "0000000000000000",
64307 => "0000000000000000",64308 => "0000000000000000",
64309 => "0000000000000000",64310 => "0000000000000000",
64311 => "0000000000000000",64312 => "0000000000000000",
64313 => "0000000000000000",64314 => "0000000000000000",
64315 => "0000000000000000",64316 => "0000000000000000",
64317 => "0000000000000000",64318 => "0000000000000000",
64319 => "0000000000000000",64320 => "0000000000000000",
64321 => "0000000000000000",64322 => "0000000000000000",
64323 => "0000000000000000",64324 => "0000000000000000",
64325 => "0000000000000000",64326 => "0000000000000000",
64327 => "0000000000000000",64328 => "0000000000000000",
64329 => "0000000000000000",64330 => "0000000000000000",
64331 => "0000000000000000",64332 => "0000000000000000",
64333 => "0000000000000000",64334 => "0000000000000000",
64335 => "0000000000000000",64336 => "0000000000000000",
64337 => "0000000000000000",64338 => "0000000000000000",
64339 => "0000000000000000",64340 => "0000000000000000",
64341 => "0000000000000000",64342 => "0000000000000000",
64343 => "0000000000000000",64344 => "0000000000000000",
64345 => "0000000000000000",64346 => "0000000000000000",
64347 => "0000000000000000",64348 => "0000000000000000",
64349 => "0000000000000000",64350 => "0000000000000000",
64351 => "0000000000000000",64352 => "0000000000000000",
64353 => "0000000000000000",64354 => "0000000000000000",
64355 => "0000000000000000",64356 => "0000000000000000",
64357 => "0000000000000000",64358 => "0000000000000000",
64359 => "0000000000000000",64360 => "0000000000000000",
64361 => "0000000000000000",64362 => "0000000000000000",
64363 => "0000000000000000",64364 => "0000000000000000",
64365 => "0000000000000000",64366 => "0000000000000000",
64367 => "0000000000000000",64368 => "0000000000000000",
64369 => "0000000000000000",64370 => "0000000000000000",
64371 => "0000000000000000",64372 => "0000000000000000",
64373 => "0000000000000000",64374 => "0000000000000000",
64375 => "0000000000000000",64376 => "0000000000000000",
64377 => "0000000000000000",64378 => "0000000000000000",
64379 => "0000000000000000",64380 => "0000000000000000",
64381 => "0000000000000000",64382 => "0000000000000000",
64383 => "0000000000000000",64384 => "0000000000000000",
64385 => "0000000000000000",64386 => "0000000000000000",
64387 => "0000000000000000",64388 => "0000000000000000",
64389 => "0000000000000000",64390 => "0000000000000000",
64391 => "0000000000000000",64392 => "0000000000000000",
64393 => "0000000000000000",64394 => "0000000000000000",
64395 => "0000000000000000",64396 => "0000000000000000",
64397 => "0000000000000000",64398 => "0000000000000000",
64399 => "0000000000000000",64400 => "0000000000000000",
64401 => "0000000000000000",64402 => "0000000000000000",
64403 => "0000000000000000",64404 => "0000000000000000",
64405 => "0000000000000000",64406 => "0000000000000000",
64407 => "0000000000000000",64408 => "0000000000000000",
64409 => "0000000000000000",64410 => "0000000000000000",
64411 => "0000000000000000",64412 => "0000000000000000",
64413 => "0000000000000000",64414 => "0000000000000000",
64415 => "0000000000000000",64416 => "0000000000000000",
64417 => "0000000000000000",64418 => "0000000000000000",
64419 => "0000000000000000",64420 => "0000000000000000",
64421 => "0000000000000000",64422 => "0000000000000000",
64423 => "0000000000000000",64424 => "0000000000000000",
64425 => "0000000000000000",64426 => "0000000000000000",
64427 => "0000000000000000",64428 => "0000000000000000",
64429 => "0000000000000000",64430 => "0000000000000000",
64431 => "0000000000000000",64432 => "0000000000000000",
64433 => "0000000000000000",64434 => "0000000000000000",
64435 => "0000000000000000",64436 => "0000000000000000",
64437 => "0000000000000000",64438 => "0000000000000000",
64439 => "0000000000000000",64440 => "0000000000000000",
64441 => "0000000000000000",64442 => "0000000000000000",
64443 => "0000000000000000",64444 => "0000000000000000",
64445 => "0000000000000000",64446 => "0000000000000000",
64447 => "0000000000000000",64448 => "0000000000000000",
64449 => "0000000000000000",64450 => "0000000000000000",
64451 => "0000000000000000",64452 => "0000000000000000",
64453 => "0000000000000000",64454 => "0000000000000000",
64455 => "0000000000000000",64456 => "0000000000000000",
64457 => "0000000000000000",64458 => "0000000000000000",
64459 => "0000000000000000",64460 => "0000000000000000",
64461 => "0000000000000000",64462 => "0000000000000000",
64463 => "0000000000000000",64464 => "0000000000000000",
64465 => "0000000000000000",64466 => "0000000000000000",
64467 => "0000000000000000",64468 => "0000000000000000",
64469 => "0000000000000000",64470 => "0000000000000000",
64471 => "0000000000000000",64472 => "0000000000000000",
64473 => "0000000000000000",64474 => "0000000000000000",
64475 => "0000000000000000",64476 => "0000000000000000",
64477 => "0000000000000000",64478 => "0000000000000000",
64479 => "0000000000000000",64480 => "0000000000000000",
64481 => "0000000000000000",64482 => "0000000000000000",
64483 => "0000000000000000",64484 => "0000000000000000",
64485 => "0000000000000000",64486 => "0000000000000000",
64487 => "0000000000000000",64488 => "0000000000000000",
64489 => "0000000000000000",64490 => "0000000000000000",
64491 => "0000000000000000",64492 => "0000000000000000",
64493 => "0000000000000000",64494 => "0000000000000000",
64495 => "0000000000000000",64496 => "0000000000000000",
64497 => "0000000000000000",64498 => "0000000000000000",
64499 => "0000000000000000",64500 => "0000000000000000",
64501 => "0000000000000000",64502 => "0000000000000000",
64503 => "0000000000000000",64504 => "0000000000000000",
64505 => "0000000000000000",64506 => "0000000000000000",
64507 => "0000000000000000",64508 => "0000000000000000",
64509 => "0000000000000000",64510 => "0000000000000000",
64511 => "0000000000000000",64512 => "0000000000000000",
64513 => "0000000000000000",64514 => "0000000000000000",
64515 => "0000000000000000",64516 => "0000000000000000",
64517 => "0000000000000000",64518 => "0000000000000000",
64519 => "0000000000000000",64520 => "0000000000000000",
64521 => "0000000000000000",64522 => "0000000000000000",
64523 => "0000000000000000",64524 => "0000000000000000",
64525 => "0000000000000000",64526 => "0000000000000000",
64527 => "0000000000000000",64528 => "0000000000000000",
64529 => "0000000000000000",64530 => "0000000000000000",
64531 => "0000000000000000",64532 => "0000000000000000",
64533 => "0000000000000000",64534 => "0000000000000000",
64535 => "0000000000000000",64536 => "0000000000000000",
64537 => "0000000000000000",64538 => "0000000000000000",
64539 => "0000000000000000",64540 => "0000000000000000",
64541 => "0000000000000000",64542 => "0000000000000000",
64543 => "0000000000000000",64544 => "0000000000000000",
64545 => "0000000000000000",64546 => "0000000000000000",
64547 => "0000000000000000",64548 => "0000000000000000",
64549 => "0000000000000000",64550 => "0000000000000000",
64551 => "0000000000000000",64552 => "0000000000000000",
64553 => "0000000000000000",64554 => "0000000000000000",
64555 => "0000000000000000",64556 => "0000000000000000",
64557 => "0000000000000000",64558 => "0000000000000000",
64559 => "0000000000000000",64560 => "0000000000000000",
64561 => "0000000000000000",64562 => "0000000000000000",
64563 => "0000000000000000",64564 => "0000000000000000",
64565 => "0000000000000000",64566 => "0000000000000000",
64567 => "0000000000000000",64568 => "0000000000000000",
64569 => "0000000000000000",64570 => "0000000000000000",
64571 => "0000000000000000",64572 => "0000000000000000",
64573 => "0000000000000000",64574 => "0000000000000000",
64575 => "0000000000000000",64576 => "0000000000000000",
64577 => "0000000000000000",64578 => "0000000000000000",
64579 => "0000000000000000",64580 => "0000000000000000",
64581 => "0000000000000000",64582 => "0000000000000000",
64583 => "0000000000000000",64584 => "0000000000000000",
64585 => "0000000000000000",64586 => "0000000000000000",
64587 => "0000000000000000",64588 => "0000000000000000",
64589 => "0000000000000000",64590 => "0000000000000000",
64591 => "0000000000000000",64592 => "0000000000000000",
64593 => "0000000000000000",64594 => "0000000000000000",
64595 => "0000000000000000",64596 => "0000000000000000",
64597 => "0000000000000000",64598 => "0000000000000000",
64599 => "0000000000000000",64600 => "0000000000000000",
64601 => "0000000000000000",64602 => "0000000000000000",
64603 => "0000000000000000",64604 => "0000000000000000",
64605 => "0000000000000000",64606 => "0000000000000000",
64607 => "0000000000000000",64608 => "0000000000000000",
64609 => "0000000000000000",64610 => "0000000000000000",
64611 => "0000000000000000",64612 => "0000000000000000",
64613 => "0000000000000000",64614 => "0000000000000000",
64615 => "0000000000000000",64616 => "0000000000000000",
64617 => "0000000000000000",64618 => "0000000000000000",
64619 => "0000000000000000",64620 => "0000000000000000",
64621 => "0000000000000000",64622 => "0000000000000000",
64623 => "0000000000000000",64624 => "0000000000000000",
64625 => "0000000000000000",64626 => "0000000000000000",
64627 => "0000000000000000",64628 => "0000000000000000",
64629 => "0000000000000000",64630 => "0000000000000000",
64631 => "0000000000000000",64632 => "0000000000000000",
64633 => "0000000000000000",64634 => "0000000000000000",
64635 => "0000000000000000",64636 => "0000000000000000",
64637 => "0000000000000000",64638 => "0000000000000000",
64639 => "0000000000000000",64640 => "0000000000000000",
64641 => "0000000000000000",64642 => "0000000000000000",
64643 => "0000000000000000",64644 => "0000000000000000",
64645 => "0000000000000000",64646 => "0000000000000000",
64647 => "0000000000000000",64648 => "0000000000000000",
64649 => "0000000000000000",64650 => "0000000000000000",
64651 => "0000000000000000",64652 => "0000000000000000",
64653 => "0000000000000000",64654 => "0000000000000000",
64655 => "0000000000000000",64656 => "0000000000000000",
64657 => "0000000000000000",64658 => "0000000000000000",
64659 => "0000000000000000",64660 => "0000000000000000",
64661 => "0000000000000000",64662 => "0000000000000000",
64663 => "0000000000000000",64664 => "0000000000000000",
64665 => "0000000000000000",64666 => "0000000000000000",
64667 => "0000000000000000",64668 => "0000000000000000",
64669 => "0000000000000000",64670 => "0000000000000000",
64671 => "0000000000000000",64672 => "0000000000000000",
64673 => "0000000000000000",64674 => "0000000000000000",
64675 => "0000000000000000",64676 => "0000000000000000",
64677 => "0000000000000000",64678 => "0000000000000000",
64679 => "0000000000000000",64680 => "0000000000000000",
64681 => "0000000000000000",64682 => "0000000000000000",
64683 => "0000000000000000",64684 => "0000000000000000",
64685 => "0000000000000000",64686 => "0000000000000000",
64687 => "0000000000000000",64688 => "0000000000000000",
64689 => "0000000000000000",64690 => "0000000000000000",
64691 => "0000000000000000",64692 => "0000000000000000",
64693 => "0000000000000000",64694 => "0000000000000000",
64695 => "0000000000000000",64696 => "0000000000000000",
64697 => "0000000000000000",64698 => "0000000000000000",
64699 => "0000000000000000",64700 => "0000000000000000",
64701 => "0000000000000000",64702 => "0000000000000000",
64703 => "0000000000000000",64704 => "0000000000000000",
64705 => "0000000000000000",64706 => "0000000000000000",
64707 => "0000000000000000",64708 => "0000000000000000",
64709 => "0000000000000000",64710 => "0000000000000000",
64711 => "0000000000000000",64712 => "0000000000000000",
64713 => "0000000000000000",64714 => "0000000000000000",
64715 => "0000000000000000",64716 => "0000000000000000",
64717 => "0000000000000000",64718 => "0000000000000000",
64719 => "0000000000000000",64720 => "0000000000000000",
64721 => "0000000000000000",64722 => "0000000000000000",
64723 => "0000000000000000",64724 => "0000000000000000",
64725 => "0000000000000000",64726 => "0000000000000000",
64727 => "0000000000000000",64728 => "0000000000000000",
64729 => "0000000000000000",64730 => "0000000000000000",
64731 => "0000000000000000",64732 => "0000000000000000",
64733 => "0000000000000000",64734 => "0000000000000000",
64735 => "0000000000000000",64736 => "0000000000000000",
64737 => "0000000000000000",64738 => "0000000000000000",
64739 => "0000000000000000",64740 => "0000000000000000",
64741 => "0000000000000000",64742 => "0000000000000000",
64743 => "0000000000000000",64744 => "0000000000000000",
64745 => "0000000000000000",64746 => "0000000000000000",
64747 => "0000000000000000",64748 => "0000000000000000",
64749 => "0000000000000000",64750 => "0000000000000000",
64751 => "0000000000000000",64752 => "0000000000000000",
64753 => "0000000000000000",64754 => "0000000000000000",
64755 => "0000000000000000",64756 => "0000000000000000",
64757 => "0000000000000000",64758 => "0000000000000000",
64759 => "0000000000000000",64760 => "0000000000000000",
64761 => "0000000000000000",64762 => "0000000000000000",
64763 => "0000000000000000",64764 => "0000000000000000",
64765 => "0000000000000000",64766 => "0000000000000000",
64767 => "0000000000000000",64768 => "0000000000000000",
64769 => "0000000000000000",64770 => "0000000000000000",
64771 => "0000000000000000",64772 => "0000000000000000",
64773 => "0000000000000000",64774 => "0000000000000000",
64775 => "0000000000000000",64776 => "0000000000000000",
64777 => "0000000000000000",64778 => "0000000000000000",
64779 => "0000000000000000",64780 => "0000000000000000",
64781 => "0000000000000000",64782 => "0000000000000000",
64783 => "0000000000000000",64784 => "0000000000000000",
64785 => "0000000000000000",64786 => "0000000000000000",
64787 => "0000000000000000",64788 => "0000000000000000",
64789 => "0000000000000000",64790 => "0000000000000000",
64791 => "0000000000000000",64792 => "0000000000000000",
64793 => "0000000000000000",64794 => "0000000000000000",
64795 => "0000000000000000",64796 => "0000000000000000",
64797 => "0000000000000000",64798 => "0000000000000000",
64799 => "0000000000000000",64800 => "0000000000000000",
64801 => "0000000000000000",64802 => "0000000000000000",
64803 => "0000000000000000",64804 => "0000000000000000",
64805 => "0000000000000000",64806 => "0000000000000000",
64807 => "0000000000000000",64808 => "0000000000000000",
64809 => "0000000000000000",64810 => "0000000000000000",
64811 => "0000000000000000",64812 => "0000000000000000",
64813 => "0000000000000000",64814 => "0000000000000000",
64815 => "0000000000000000",64816 => "0000000000000000",
64817 => "0000000000000000",64818 => "0000000000000000",
64819 => "0000000000000000",64820 => "0000000000000000",
64821 => "0000000000000000",64822 => "0000000000000000",
64823 => "0000000000000000",64824 => "0000000000000000",
64825 => "0000000000000000",64826 => "0000000000000000",
64827 => "0000000000000000",64828 => "0000000000000000",
64829 => "0000000000000000",64830 => "0000000000000000",
64831 => "0000000000000000",64832 => "0000000000000000",
64833 => "0000000000000000",64834 => "0000000000000000",
64835 => "0000000000000000",64836 => "0000000000000000",
64837 => "0000000000000000",64838 => "0000000000000000",
64839 => "0000000000000000",64840 => "0000000000000000",
64841 => "0000000000000000",64842 => "0000000000000000",
64843 => "0000000000000000",64844 => "0000000000000000",
64845 => "0000000000000000",64846 => "0000000000000000",
64847 => "0000000000000000",64848 => "0000000000000000",
64849 => "0000000000000000",64850 => "0000000000000000",
64851 => "0000000000000000",64852 => "0000000000000000",
64853 => "0000000000000000",64854 => "0000000000000000",
64855 => "0000000000000000",64856 => "0000000000000000",
64857 => "0000000000000000",64858 => "0000000000000000",
64859 => "0000000000000000",64860 => "0000000000000000",
64861 => "0000000000000000",64862 => "0000000000000000",
64863 => "0000000000000000",64864 => "0000000000000000",
64865 => "0000000000000000",64866 => "0000000000000000",
64867 => "0000000000000000",64868 => "0000000000000000",
64869 => "0000000000000000",64870 => "0000000000000000",
64871 => "0000000000000000",64872 => "0000000000000000",
64873 => "0000000000000000",64874 => "0000000000000000",
64875 => "0000000000000000",64876 => "0000000000000000",
64877 => "0000000000000000",64878 => "0000000000000000",
64879 => "0000000000000000",64880 => "0000000000000000",
64881 => "0000000000000000",64882 => "0000000000000000",
64883 => "0000000000000000",64884 => "0000000000000000",
64885 => "0000000000000000",64886 => "0000000000000000",
64887 => "0000000000000000",64888 => "0000000000000000",
64889 => "0000000000000000",64890 => "0000000000000000",
64891 => "0000000000000000",64892 => "0000000000000000",
64893 => "0000000000000000",64894 => "0000000000000000",
64895 => "0000000000000000",64896 => "0000000000000000",
64897 => "0000000000000000",64898 => "0000000000000000",
64899 => "0000000000000000",64900 => "0000000000000000",
64901 => "0000000000000000",64902 => "0000000000000000",
64903 => "0000000000000000",64904 => "0000000000000000",
64905 => "0000000000000000",64906 => "0000000000000000",
64907 => "0000000000000000",64908 => "0000000000000000",
64909 => "0000000000000000",64910 => "0000000000000000",
64911 => "0000000000000000",64912 => "0000000000000000",
64913 => "0000000000000000",64914 => "0000000000000000",
64915 => "0000000000000000",64916 => "0000000000000000",
64917 => "0000000000000000",64918 => "0000000000000000",
64919 => "0000000000000000",64920 => "0000000000000000",
64921 => "0000000000000000",64922 => "0000000000000000",
64923 => "0000000000000000",64924 => "0000000000000000",
64925 => "0000000000000000",64926 => "0000000000000000",
64927 => "0000000000000000",64928 => "0000000000000000",
64929 => "0000000000000000",64930 => "0000000000000000",
64931 => "0000000000000000",64932 => "0000000000000000",
64933 => "0000000000000000",64934 => "0000000000000000",
64935 => "0000000000000000",64936 => "0000000000000000",
64937 => "0000000000000000",64938 => "0000000000000000",
64939 => "0000000000000000",64940 => "0000000000000000",
64941 => "0000000000000000",64942 => "0000000000000000",
64943 => "0000000000000000",64944 => "0000000000000000",
64945 => "0000000000000000",64946 => "0000000000000000",
64947 => "0000000000000000",64948 => "0000000000000000",
64949 => "0000000000000000",64950 => "0000000000000000",
64951 => "0000000000000000",64952 => "0000000000000000",
64953 => "0000000000000000",64954 => "0000000000000000",
64955 => "0000000000000000",64956 => "0000000000000000",
64957 => "0000000000000000",64958 => "0000000000000000",
64959 => "0000000000000000",64960 => "0000000000000000",
64961 => "0000000000000000",64962 => "0000000000000000",
64963 => "0000000000000000",64964 => "0000000000000000",
64965 => "0000000000000000",64966 => "0000000000000000",
64967 => "0000000000000000",64968 => "0000000000000000",
64969 => "0000000000000000",64970 => "0000000000000000",
64971 => "0000000000000000",64972 => "0000000000000000",
64973 => "0000000000000000",64974 => "0000000000000000",
64975 => "0000000000000000",64976 => "0000000000000000",
64977 => "0000000000000000",64978 => "0000000000000000",
64979 => "0000000000000000",64980 => "0000000000000000",
64981 => "0000000000000000",64982 => "0000000000000000",
64983 => "0000000000000000",64984 => "0000000000000000",
64985 => "0000000000000000",64986 => "0000000000000000",
64987 => "0000000000000000",64988 => "0000000000000000",
64989 => "0000000000000000",64990 => "0000000000000000",
64991 => "0000000000000000",64992 => "0000000000000000",
64993 => "0000000000000000",64994 => "0000000000000000",
64995 => "0000000000000000",64996 => "0000000000000000",
64997 => "0000000000000000",64998 => "0000000000000000",
64999 => "0000000000000000",65000 => "0000000000000000",
65001 => "0000000000000000",65002 => "0000000000000000",
65003 => "0000000000000000",65004 => "0000000000000000",
65005 => "0000000000000000",65006 => "0000000000000000",
65007 => "0000000000000000",65008 => "0000000000000000",
65009 => "0000000000000000",65010 => "0000000000000000",
65011 => "0000000000000000",65012 => "0000000000000000",
65013 => "0000000000000000",65014 => "0000000000000000",
65015 => "0000000000000000",65016 => "0000000000000000",
65017 => "0000000000000000",65018 => "0000000000000000",
65019 => "0000000000000000",65020 => "0000000000000000",
65021 => "0000000000000000",65022 => "0000000000000000",
65023 => "0000000000000000",65024 => "0000000000000000",
65025 => "0000000000000000",65026 => "0000000000000000",
65027 => "0000000000000000",65028 => "0000000000000000",
65029 => "0000000000000000",65030 => "0000000000000000",
65031 => "0000000000000000",65032 => "0000000000000000",
65033 => "0000000000000000",65034 => "0000000000000000",
65035 => "0000000000000000",65036 => "0000000000000000",
65037 => "0000000000000000",65038 => "0000000000000000",
65039 => "0000000000000000",65040 => "0000000000000000",
65041 => "0000000000000000",65042 => "0000000000000000",
65043 => "0000000000000000",65044 => "0000000000000000",
65045 => "0000000000000000",65046 => "0000000000000000",
65047 => "0000000000000000",65048 => "0000000000000000",
65049 => "0000000000000000",65050 => "0000000000000000",
65051 => "0000000000000000",65052 => "0000000000000000",
65053 => "0000000000000000",65054 => "0000000000000000",
65055 => "0000000000000000",65056 => "0000000000000000",
65057 => "0000000000000000",65058 => "0000000000000000",
65059 => "0000000000000000",65060 => "0000000000000000",
65061 => "0000000000000000",65062 => "0000000000000000",
65063 => "0000000000000000",65064 => "0000000000000000",
65065 => "0000000000000000",65066 => "0000000000000000",
65067 => "0000000000000000",65068 => "0000000000000000",
65069 => "0000000000000000",65070 => "0000000000000000",
65071 => "0000000000000000",65072 => "0000000000000000",
65073 => "0000000000000000",65074 => "0000000000000000",
65075 => "0000000000000000",65076 => "0000000000000000",
65077 => "0000000000000000",65078 => "0000000000000000",
65079 => "0000000000000000",65080 => "0000000000000000",
65081 => "0000000000000000",65082 => "0000000000000000",
65083 => "0000000000000000",65084 => "0000000000000000",
65085 => "0000000000000000",65086 => "0000000000000000",
65087 => "0000000000000000",65088 => "0000000000000000",
65089 => "0000000000000000",65090 => "0000000000000000",
65091 => "0000000000000000",65092 => "0000000000000000",
65093 => "0000000000000000",65094 => "0000000000000000",
65095 => "0000000000000000",65096 => "0000000000000000",
65097 => "0000000000000000",65098 => "0000000000000000",
65099 => "0000000000000000",65100 => "0000000000000000",
65101 => "0000000000000000",65102 => "0000000000000000",
65103 => "0000000000000000",65104 => "0000000000000000",
65105 => "0000000000000000",65106 => "0000000000000000",
65107 => "0000000000000000",65108 => "0000000000000000",
65109 => "0000000000000000",65110 => "0000000000000000",
65111 => "0000000000000000",65112 => "0000000000000000",
65113 => "0000000000000000",65114 => "0000000000000000",
65115 => "0000000000000000",65116 => "0000000000000000",
65117 => "0000000000000000",65118 => "0000000000000000",
65119 => "0000000000000000",65120 => "0000000000000000",
65121 => "0000000000000000",65122 => "0000000000000000",
65123 => "0000000000000000",65124 => "0000000000000000",
65125 => "0000000000000000",65126 => "0000000000000000",
65127 => "0000000000000000",65128 => "0000000000000000",
65129 => "0000000000000000",65130 => "0000000000000000",
65131 => "0000000000000000",65132 => "0000000000000000",
65133 => "0000000000000000",65134 => "0000000000000000",
65135 => "0000000000000000",65136 => "0000000000000000",
65137 => "0000000000000000",65138 => "0000000000000000",
65139 => "0000000000000000",65140 => "0000000000000000",
65141 => "0000000000000000",65142 => "0000000000000000",
65143 => "0000000000000000",65144 => "0000000000000000",
65145 => "0000000000000000",65146 => "0000000000000000",
65147 => "0000000000000000",65148 => "0000000000000000",
65149 => "0000000000000000",65150 => "0000000000000000",
65151 => "0000000000000000",65152 => "0000000000000000",
65153 => "0000000000000000",65154 => "0000000000000000",
65155 => "0000000000000000",65156 => "0000000000000000",
65157 => "0000000000000000",65158 => "0000000000000000",
65159 => "0000000000000000",65160 => "0000000000000000",
65161 => "0000000000000000",65162 => "0000000000000000",
65163 => "0000000000000000",65164 => "0000000000000000",
65165 => "0000000000000000",65166 => "0000000000000000",
65167 => "0000000000000000",65168 => "0000000000000000",
65169 => "0000000000000000",65170 => "0000000000000000",
65171 => "0000000000000000",65172 => "0000000000000000",
65173 => "0000000000000000",65174 => "0000000000000000",
65175 => "0000000000000000",65176 => "0000000000000000",
65177 => "0000000000000000",65178 => "0000000000000000",
65179 => "0000000000000000",65180 => "0000000000000000",
65181 => "0000000000000000",65182 => "0000000000000000",
65183 => "0000000000000000",65184 => "0000000000000000",
65185 => "0000000000000000",65186 => "0000000000000000",
65187 => "0000000000000000",65188 => "0000000000000000",
65189 => "0000000000000000",65190 => "0000000000000000",
65191 => "0000000000000000",65192 => "0000000000000000",
65193 => "0000000000000000",65194 => "0000000000000000",
65195 => "0000000000000000",65196 => "0000000000000000",
65197 => "0000000000000000",65198 => "0000000000000000",
65199 => "0000000000000000",65200 => "0000000000000000",
65201 => "0000000000000000",65202 => "0000000000000000",
65203 => "0000000000000000",65204 => "0000000000000000",
65205 => "0000000000000000",65206 => "0000000000000000",
65207 => "0000000000000000",65208 => "0000000000000000",
65209 => "0000000000000000",65210 => "0000000000000000",
65211 => "0000000000000000",65212 => "0000000000000000",
65213 => "0000000000000000",65214 => "0000000000000000",
65215 => "0000000000000000",65216 => "0000000000000000",
65217 => "0000000000000000",65218 => "0000000000000000",
65219 => "0000000000000000",65220 => "0000000000000000",
65221 => "0000000000000000",65222 => "0000000000000000",
65223 => "0000000000000000",65224 => "0000000000000000",
65225 => "0000000000000000",65226 => "0000000000000000",
65227 => "0000000000000000",65228 => "0000000000000000",
65229 => "0000000000000000",65230 => "0000000000000000",
65231 => "0000000000000000",65232 => "0000000000000000",
65233 => "0000000000000000",65234 => "0000000000000000",
65235 => "0000000000000000",65236 => "0000000000000000",
65237 => "0000000000000000",65238 => "0000000000000000",
65239 => "0000000000000000",65240 => "0000000000000000",
65241 => "0000000000000000",65242 => "0000000000000000",
65243 => "0000000000000000",65244 => "0000000000000000",
65245 => "0000000000000000",65246 => "0000000000000000",
65247 => "0000000000000000",65248 => "0000000000000000",
65249 => "0000000000000000",65250 => "0000000000000000",
65251 => "0000000000000000",65252 => "0000000000000000",
65253 => "0000000000000000",65254 => "0000000000000000",
65255 => "0000000000000000",65256 => "0000000000000000",
65257 => "0000000000000000",65258 => "0000000000000000",
65259 => "0000000000000000",65260 => "0000000000000000",
65261 => "0000000000000000",65262 => "0000000000000000",
65263 => "0000000000000000",65264 => "0000000000000000",
65265 => "0000000000000000",65266 => "0000000000000000",
65267 => "0000000000000000",65268 => "0000000000000000",
65269 => "0000000000000000",65270 => "0000000000000000",
65271 => "0000000000000000",65272 => "0000000000000000",
65273 => "0000000000000000",65274 => "0000000000000000",
65275 => "0000000000000000",65276 => "0000000000000000",
65277 => "0000000000000000",65278 => "0000000000000000",
65279 => "0000000000000000",65280 => "0000000000000000",
65281 => "0000000000000000",65282 => "0000000000000000",
65283 => "0000000000000000",65284 => "0000000000000000",
65285 => "0000000000000000",65286 => "0000000000000000",
65287 => "0000000000000000",65288 => "0000000000000000",
65289 => "0000000000000000",65290 => "0000000000000000",
65291 => "0000000000000000",65292 => "0000000000000000",
65293 => "0000000000000000",65294 => "0000000000000000",
65295 => "0000000000000000",65296 => "0000000000000000",
65297 => "0000000000000000",65298 => "0000000000000000",
65299 => "0000000000000000",65300 => "0000000000000000",
65301 => "0000000000000000",65302 => "0000000000000000",
65303 => "0000000000000000",65304 => "0000000000000000",
65305 => "0000000000000000",65306 => "0000000000000000",
65307 => "0000000000000000",65308 => "0000000000000000",
65309 => "0000000000000000",65310 => "0000000000000000",
65311 => "0000000000000000",65312 => "0000000000000000",
65313 => "0000000000000000",65314 => "0000000000000000",
65315 => "0000000000000000",65316 => "0000000000000000",
65317 => "0000000000000000",65318 => "0000000000000000",
65319 => "0000000000000000",65320 => "0000000000000000",
65321 => "0000000000000000",65322 => "0000000000000000",
65323 => "0000000000000000",65324 => "0000000000000000",
65325 => "0000000000000000",65326 => "0000000000000000",
65327 => "0000000000000000",65328 => "0000000000000000",
65329 => "0000000000000000",65330 => "0000000000000000",
65331 => "0000000000000000",65332 => "0000000000000000",
65333 => "0000000000000000",65334 => "0000000000000000",
65335 => "0000000000000000",65336 => "0000000000000000",
65337 => "0000000000000000",65338 => "0000000000000000",
65339 => "0000000000000000",65340 => "0000000000000000",
65341 => "0000000000000000",65342 => "0000000000000000",
65343 => "0000000000000000",65344 => "0000000000000000",
65345 => "0000000000000000",65346 => "0000000000000000",
65347 => "0000000000000000",65348 => "0000000000000000",
65349 => "0000000000000000",65350 => "0000000000000000",
65351 => "0000000000000000",65352 => "0000000000000000",
65353 => "0000000000000000",65354 => "0000000000000000",
65355 => "0000000000000000",65356 => "0000000000000000",
65357 => "0000000000000000",65358 => "0000000000000000",
65359 => "0000000000000000",65360 => "0000000000000000",
65361 => "0000000000000000",65362 => "0000000000000000",
65363 => "0000000000000000",65364 => "0000000000000000",
65365 => "0000000000000000",65366 => "0000000000000000",
65367 => "0000000000000000",65368 => "0000000000000000",
65369 => "0000000000000000",65370 => "0000000000000000",
65371 => "0000000000000000",65372 => "0000000000000000",
65373 => "0000000000000000",65374 => "0000000000000000",
65375 => "0000000000000000",65376 => "0000000000000000",
65377 => "0000000000000000",65378 => "0000000000000000",
65379 => "0000000000000000",65380 => "0000000000000000",
65381 => "0000000000000000",65382 => "0000000000000000",
65383 => "0000000000000000",65384 => "0000000000000000",
65385 => "0000000000000000",65386 => "0000000000000000",
65387 => "0000000000000000",65388 => "0000000000000000",
65389 => "0000000000000000",65390 => "0000000000000000",
65391 => "0000000000000000",65392 => "0000000000000000",
65393 => "0000000000000000",65394 => "0000000000000000",
65395 => "0000000000000000",65396 => "0000000000000000",
65397 => "0000000000000000",65398 => "0000000000000000",
65399 => "0000000000000000",65400 => "0000000000000000",
65401 => "0000000000000000",65402 => "0000000000000000",
65403 => "0000000000000000",65404 => "0000000000000000",
65405 => "0000000000000000",65406 => "0000000000000000",
65407 => "0000000000000000",65408 => "0000000000000000",
65409 => "0000000000000000",65410 => "0000000000000000",
65411 => "0000000000000000",65412 => "0000000000000000",
65413 => "0000000000000000",65414 => "0000000000000000",
65415 => "0000000000000000",65416 => "0000000000000000",
65417 => "0000000000000000",65418 => "0000000000000000",
65419 => "0000000000000000",65420 => "0000000000000000",
65421 => "0000000000000000",65422 => "0000000000000000",
65423 => "0000000000000000",65424 => "0000000000000000",
65425 => "0000000000000000",65426 => "0000000000000000",
65427 => "0000000000000000",65428 => "0000000000000000",
65429 => "0000000000000000",65430 => "0000000000000000",
65431 => "0000000000000000",65432 => "0000000000000000",
65433 => "0000000000000000",65434 => "0000000000000000",
65435 => "0000000000000000",65436 => "0000000000000000",
65437 => "0000000000000000",65438 => "0000000000000000",
65439 => "0000000000000000",65440 => "0000000000000000",
65441 => "0000000000000000",65442 => "0000000000000000",
65443 => "0000000000000000",65444 => "0000000000000000",
65445 => "0000000000000000",65446 => "0000000000000000",
65447 => "0000000000000000",65448 => "0000000000000000",
65449 => "0000000000000000",65450 => "0000000000000000",
65451 => "0000000000000000",65452 => "0000000000000000",
65453 => "0000000000000000",65454 => "0000000000000000",
65455 => "0000000000000000",65456 => "0000000000000000",
65457 => "0000000000000000",65458 => "0000000000000000",
65459 => "0000000000000000",65460 => "0000000000000000",
65461 => "0000000000000000",65462 => "0000000000000000",
65463 => "0000000000000000",65464 => "0000000000000000",
65465 => "0000000000000000",65466 => "0000000000000000",
65467 => "0000000000000000",65468 => "0000000000000000",
65469 => "0000000000000000",65470 => "0000000000000000",
65471 => "0000000000000000",65472 => "0000000000000000",
65473 => "0000000000000000",65474 => "0000000000000000",
65475 => "0000000000000000",65476 => "0000000000000000",
65477 => "0000000000000000",65478 => "0000000000000000",
65479 => "0000000000000000",65480 => "0000000000000000",
65481 => "0000000000000000",65482 => "0000000000000000",
65483 => "0000000000000000",65484 => "0000000000000000",
65485 => "0000000000000000",65486 => "0000000000000000",
65487 => "0000000000000000",65488 => "0000000000000000",
65489 => "0000000000000000",65490 => "0000000000000000",
65491 => "0000000000000000",65492 => "0000000000000000",
65493 => "0000000000000000",65494 => "0000000000000000",
65495 => "0000000000000000",65496 => "0000000000000000",
65497 => "0000000000000000",65498 => "0000000000000000",
65499 => "0000000000000000",65500 => "0000000000000000",
65501 => "0000000000000000",65502 => "0000000000000000",
65503 => "0000000000000000",65504 => "0000000000000000",
65505 => "0000000000000000",65506 => "0000000000000000",
65507 => "0000000000000000",65508 => "0000000000000000",
65509 => "0000000000000000",65510 => "0000000000000000",
65511 => "0000000000000000",65512 => "0000000000000000",
65513 => "0000000000000000",65514 => "0000000000000000",
65515 => "0000000000000000",65516 => "0000000000000000",
65517 => "0000000000000000",65518 => "0000000000000000",
65519 => "0000000000000000",65520 => "0000000000000000",
65521 => "0000000000000000",65522 => "0000000000000000",
65523 => "0000000000000000",65524 => "0000000000000000",
65525 => "0000000000000000",65526 => "0000000000000000",
65527 => "0000000000000000",65528 => "0000000000000000",
65529 => "0000000000000000",65530 => "0000000000000000",
65531 => "0000000000000000",65532 => "0000000000000000",
65533 => "0000000000000000",65534 => "0000000000000000",
65535 => "0000000000000000");
begin

	findValue: process (clk,bitVector) is 
		variable index : integer := 0;

		BEGIN  
			index := to_integer(unsigned(bitVector));
			outVector <= exp_lut(index);

	end process findValue;

end architecture;

