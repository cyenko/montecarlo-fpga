----------------------------------------------------------------------------- 
library IEEE; 
 
use IEEE.std_logic_1164.all; 
use WORK.monte_carlo.all; 
--Additional standard or custom libraries go here 
use IEEE.numeric_std.all;

--inputs: clock, start, stock price, strike, t
--output: premium, stock price out, ready
--	for now, do only premium and ready

entity exp is 
 port( 
	 --Inputs 
	 clk : in std_logic; 
	 bitVector : in std_logic_vector (15 downto 0); --16 bits
	 
	 --Outputs 
	 outVector : out std_logic_vector (15 downto 0)
 ); 
end entity exp;

architecture behavioral of exp is 
--Declare the ROM type
type rom is array (0 to 2**16-1) of std_logic_vector(15 downto 0);
--Input the LUT, this will be generated by python
constant exp_lut : rom := (0=>"0000000000000000",1=>"0000000000000001");

begin

	findValue: process (clk,bitVector) is 
		variable index : integer := 0;

		BEGIN  
			index := to_integer(bitVector);
			outVector <= exp_lut(index);

	end process findValue;

end architecture;

