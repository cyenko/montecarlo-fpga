----------------------------------------------------------------------------- 
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_unsigned.all;
use work.monte_carlo.all;

--inputs: clock, start, stock price, strike, t
--output: premium, stock price out, ready
--	for now, do only premium and ready

entity exp_fn is 
 port( 
	 --Inputs 
	 clk : in std_logic; 
	 bitVector : in std_logic_vector (15 downto 0); --16 bits
	 
	 --Outputs 
	 outVector : out std_logic_vector (15 downto 0)
 ); 
end entity exp_fn;

architecture behavioral of exp_fn is 
--Declare the ROM type
--Real length will be 0 to 2**16-1
--type rom is array (0 to (2**16)-1) of std_logic_vector(15 downto 0);
type rom is array (0 to (3414)) of std_logic_vector(15 downto 0);
type rom_n is array(32768 to 34194) of std_logic_vector(15 downto 0);
--Input the LUT, this will be generated by python
--constant exp_lut : rom := (0=>"0000000000000000",1=>"0000000000000001");
constant exp_lut : rom := (0 => "0000000100000000",
	1 => "0000000100000001",2 => "0000000100000010",3 => "0000000100000011",
	4 => "0000000100000100",5 => "0000000100000101",6 => "0000000100000110",
	7 => "0000000100000111",8 => "0000000100001000",9 => "0000000100001001",
	10 => "0000000100001010",11 => "0000000100001011",12 => "0000000100001100",
	13 => "0000000100001101",14 => "0000000100001110",15 => "0000000100001111",
	16 => "0000000100010000",17 => "0000000100010001",18 => "0000000100010010",
	19 => "0000000100010011",20 => "0000000100010100",21 => "0000000100010101",
	22 => "0000000100010110",23 => "0000000100011000",24 => "0000000100011001",
	25 => "0000000100011010",26 => "0000000100011011",27 => "0000000100011100",
	28 => "0000000100011101",29 => "0000000100011110",30 => "0000000100011111",
	31 => "0000000100100000",32 => "0000000100100010",33 => "0000000100100011",
	34 => "0000000100100100",35 => "0000000100100101",36 => "0000000100100110",
	37 => "0000000100100111",38 => "0000000100101000",39 => "0000000100101010",
	40 => "0000000100101011",41 => "0000000100101100",42 => "0000000100101101",
	43 => "0000000100101110",44 => "0000000100110000",45 => "0000000100110001",
	46 => "0000000100110010",47 => "0000000100110011",48 => "0000000100110100",
	49 => "0000000100110110",50 => "0000000100110111",51 => "0000000100111000",
	52 => "0000000100111001",53 => "0000000100111010",54 => "0000000100111100",
	55 => "0000000100111101",56 => "0000000100111110",57 => "0000000100111111",
	58 => "0000000101000001",59 => "0000000101000010",60 => "0000000101000011",
	61 => "0000000101000100",62 => "0000000101000110",63 => "0000000101000111",
	64 => "0000000101001000",65 => "0000000101001001",66 => "0000000101001011",
	67 => "0000000101001100",68 => "0000000101001101",69 => "0000000101001111",
	70 => "0000000101010000",71 => "0000000101010001",72 => "0000000101010011",
	73 => "0000000101010100",74 => "0000000101010101",75 => "0000000101010111",
	76 => "0000000101011000",77 => "0000000101011001",78 => "0000000101011011",
	79 => "0000000101011100",80 => "0000000101011101",81 => "0000000101011111",
	82 => "0000000101100000",83 => "0000000101100010",84 => "0000000101100011",
	85 => "0000000101100100",86 => "0000000101100110",87 => "0000000101100111",
	88 => "0000000101101001",89 => "0000000101101010",90 => "0000000101101011",
	91 => "0000000101101101",92 => "0000000101101110",93 => "0000000101110000",
	94 => "0000000101110001",95 => "0000000101110011",96 => "0000000101110100",
	97 => "0000000101110101",98 => "0000000101110111",99 => "0000000101111000",
	100 => "0000000101111010",101 => "0000000101111011",102 => "0000000101111101",
	103 => "0000000101111110",104 => "0000000110000000",105 => "0000000110000001",
	106 => "0000000110000011",107 => "0000000110000100",108 => "0000000110000110",
	109 => "0000000110000111",110 => "0000000110001001",111 => "0000000110001010",
	112 => "0000000110001100",113 => "0000000110001110",114 => "0000000110001111",
	115 => "0000000110010001",116 => "0000000110010010",117 => "0000000110010100",
	118 => "0000000110010101",119 => "0000000110010111",120 => "0000000110011001",
	121 => "0000000110011010",122 => "0000000110011100",123 => "0000000110011101",
	124 => "0000000110011111",125 => "0000000110100001",126 => "0000000110100010",
	127 => "0000000110100100",128 => "0000000110100110",129 => "0000000110100111",
	130 => "0000000110101001",131 => "0000000110101011",132 => "0000000110101100",
	133 => "0000000110101110",134 => "0000000110110000",135 => "0000000110110001",
	136 => "0000000110110011",137 => "0000000110110101",138 => "0000000110110110",
	139 => "0000000110111000",140 => "0000000110111010",141 => "0000000110111100",
	142 => "0000000110111101",143 => "0000000110111111",144 => "0000000111000001",
	145 => "0000000111000011",146 => "0000000111000100",147 => "0000000111000110",
	148 => "0000000111001000",149 => "0000000111001010",150 => "0000000111001011",
	151 => "0000000111001101",152 => "0000000111001111",153 => "0000000111010001",
	154 => "0000000111010011",155 => "0000000111010101",156 => "0000000111010110",
	157 => "0000000111011000",158 => "0000000111011010",159 => "0000000111011100",
	160 => "0000000111011110",161 => "0000000111100000",162 => "0000000111100010",
	163 => "0000000111100011",164 => "0000000111100101",165 => "0000000111100111",
	166 => "0000000111101001",167 => "0000000111101011",168 => "0000000111101101",
	169 => "0000000111101111",170 => "0000000111110001",171 => "0000000111110011",
	172 => "0000000111110101",173 => "0000000111110111",174 => "0000000111111001",
	175 => "0000000111111011",176 => "0000000111111101",177 => "0000000111111111",
	178 => "0000001000000001",179 => "0000001000000011",180 => "0000001000000101",
	181 => "0000001000000111",182 => "0000001000001001",183 => "0000001000001011",
	184 => "0000001000001101",185 => "0000001000001111",186 => "0000001000010001",
	187 => "0000001000010011",188 => "0000001000010101",189 => "0000001000010111",
	190 => "0000001000011001",191 => "0000001000011011",192 => "0000001000011101",
	193 => "0000001000100000",194 => "0000001000100010",195 => "0000001000100100",
	196 => "0000001000100110",197 => "0000001000101000",198 => "0000001000101010",
	199 => "0000001000101100",200 => "0000001000101111",201 => "0000001000110001",
	202 => "0000001000110011",203 => "0000001000110101",204 => "0000001000110111",
	205 => "0000001000111010",206 => "0000001000111100",207 => "0000001000111110",
	208 => "0000001001000000",209 => "0000001001000011",210 => "0000001001000101",
	211 => "0000001001000111",212 => "0000001001001001",213 => "0000001001001100",
	214 => "0000001001001110",215 => "0000001001010000",216 => "0000001001010011",
	217 => "0000001001010101",218 => "0000001001010111",219 => "0000001001011010",
	220 => "0000001001011100",221 => "0000001001011110",222 => "0000001001100001",
	223 => "0000001001100011",224 => "0000001001100110",225 => "0000001001101000",
	226 => "0000001001101010",227 => "0000001001101101",228 => "0000001001101111",
	229 => "0000001001110010",230 => "0000001001110100",231 => "0000001001110111",
	232 => "0000001001111001",233 => "0000001001111100",234 => "0000001001111110",
	235 => "0000001010000001",236 => "0000001010000011",237 => "0000001010000110",
	238 => "0000001010001000",239 => "0000001010001011",240 => "0000001010001101",
	241 => "0000001010010000",242 => "0000001010010010",243 => "0000001010010101",
	244 => "0000001010011000",245 => "0000001010011010",246 => "0000001010011101",
	247 => "0000001010011111",248 => "0000001010100010",249 => "0000001010100101",
	250 => "0000001010100111",251 => "0000001010101010",252 => "0000001010101101",
	253 => "0000001010101111",254 => "0000001010110010",255 => "0000001010110101",
	256 => "0000001010110111",257 => "0000001010111010",258 => "0000001010111101",
	259 => "0000001011000000",260 => "0000001011000010",261 => "0000001011000101",
	262 => "0000001011001000",263 => "0000001011001011",264 => "0000001011001101",
	265 => "0000001011010000",266 => "0000001011010011",267 => "0000001011010110",
	268 => "0000001011011001",269 => "0000001011011100",270 => "0000001011011110",
	271 => "0000001011100001",272 => "0000001011100100",273 => "0000001011100111",
	274 => "0000001011101010",275 => "0000001011101101",276 => "0000001011110000",
	277 => "0000001011110011",278 => "0000001011110110",279 => "0000001011111001",
	280 => "0000001011111100",281 => "0000001011111111",282 => "0000001100000010",
	283 => "0000001100000101",284 => "0000001100001000",285 => "0000001100001011",
	286 => "0000001100001110",287 => "0000001100010001",288 => "0000001100010100",
	289 => "0000001100010111",290 => "0000001100011010",291 => "0000001100011101",
	292 => "0000001100100000",293 => "0000001100100100",294 => "0000001100100111",
	295 => "0000001100101010",296 => "0000001100101101",297 => "0000001100110000",
	298 => "0000001100110011",299 => "0000001100110111",300 => "0000001100111010",
	301 => "0000001100111101",302 => "0000001101000000",303 => "0000001101000100",
	304 => "0000001101000111",305 => "0000001101001010",306 => "0000001101001101",
	307 => "0000001101010001",308 => "0000001101010100",309 => "0000001101010111",
	310 => "0000001101011011",311 => "0000001101011110",312 => "0000001101100010",
	313 => "0000001101100101",314 => "0000001101101000",315 => "0000001101101100",
	316 => "0000001101101111",317 => "0000001101110011",318 => "0000001101110110",
	319 => "0000001101111010",320 => "0000001101111101",321 => "0000001110000001",
	322 => "0000001110000100",323 => "0000001110001000",324 => "0000001110001011",
	325 => "0000001110001111",326 => "0000001110010010",327 => "0000001110010110",
	328 => "0000001110011001",329 => "0000001110011101",330 => "0000001110100001",
	331 => "0000001110100100",332 => "0000001110101000",333 => "0000001110101100",
	334 => "0000001110101111",335 => "0000001110110011",336 => "0000001110110111",
	337 => "0000001110111010",338 => "0000001110111110",339 => "0000001111000010",
	340 => "0000001111000110",341 => "0000001111001001",342 => "0000001111001101",
	343 => "0000001111010001",344 => "0000001111010101",345 => "0000001111011001",
	346 => "0000001111011101",347 => "0000001111100000",348 => "0000001111100100",
	349 => "0000001111101000",350 => "0000001111101100",351 => "0000001111110000",
	352 => "0000001111110100",353 => "0000001111111000",354 => "0000001111111100",
	355 => "0000010000000000",356 => "0000010000000100",357 => "0000010000001000",
	358 => "0000010000001100",359 => "0000010000010000",360 => "0000010000010100",
	361 => "0000010000011000",362 => "0000010000011100",363 => "0000010000100000",
	364 => "0000010000100101",365 => "0000010000101001",366 => "0000010000101101",
	367 => "0000010000110001",368 => "0000010000110101",369 => "0000010000111010",
	370 => "0000010000111110",371 => "0000010001000010",372 => "0000010001000110",
	373 => "0000010001001011",374 => "0000010001001111",375 => "0000010001010011",
	376 => "0000010001011000",377 => "0000010001011100",378 => "0000010001100000",
	379 => "0000010001100101",380 => "0000010001101001",381 => "0000010001101101",
	382 => "0000010001110010",383 => "0000010001110110",384 => "0000010001111011",
	385 => "0000010001111111",386 => "0000010010000100",387 => "0000010010001000",
	388 => "0000010010001101",389 => "0000010010010001",390 => "0000010010010110",
	391 => "0000010010011011",392 => "0000010010011111",393 => "0000010010100100",
	394 => "0000010010101001",395 => "0000010010101101",396 => "0000010010110010",
	397 => "0000010010110111",398 => "0000010010111011",399 => "0000010011000000",
	400 => "0000010011000101",401 => "0000010011001010",402 => "0000010011001110",
	403 => "0000010011010011",404 => "0000010011011000",405 => "0000010011011101",
	406 => "0000010011100010",407 => "0000010011100111",408 => "0000010011101100",
	409 => "0000010011110001",410 => "0000010011110101",411 => "0000010011111010",
	412 => "0000010011111111",413 => "0000010100000100",414 => "0000010100001001",
	415 => "0000010100001111",416 => "0000010100010100",417 => "0000010100011001",
	418 => "0000010100011110",419 => "0000010100100011",420 => "0000010100101000",
	421 => "0000010100101101",422 => "0000010100110010",423 => "0000010100111000",
	424 => "0000010100111101",425 => "0000010101000010",426 => "0000010101000111",
	427 => "0000010101001101",428 => "0000010101010010",429 => "0000010101010111",
	430 => "0000010101011101",431 => "0000010101100010",432 => "0000010101100111",
	433 => "0000010101101101",434 => "0000010101110010",435 => "0000010101111000",
	436 => "0000010101111101",437 => "0000010110000011",438 => "0000010110001000",
	439 => "0000010110001110",440 => "0000010110010011",441 => "0000010110011001",
	442 => "0000010110011111",443 => "0000010110100100",444 => "0000010110101010",
	445 => "0000010110110000",446 => "0000010110110101",447 => "0000010110111011",
	448 => "0000010111000001",449 => "0000010111000110",450 => "0000010111001100",
	451 => "0000010111010010",452 => "0000010111011000",453 => "0000010111011110",
	454 => "0000010111100100",455 => "0000010111101010",456 => "0000010111101111",
	457 => "0000010111110101",458 => "0000010111111011",459 => "0000011000000001",
	460 => "0000011000000111",461 => "0000011000001101",462 => "0000011000010011",
	463 => "0000011000011010",464 => "0000011000100000",465 => "0000011000100110",
	466 => "0000011000101100",467 => "0000011000110010",468 => "0000011000111000",
	469 => "0000011000111111",470 => "0000011001000101",471 => "0000011001001011",
	472 => "0000011001010001",473 => "0000011001011000",474 => "0000011001011110",
	475 => "0000011001100101",476 => "0000011001101011",477 => "0000011001110001",
	478 => "0000011001111000",479 => "0000011001111110",480 => "0000011010000101",
	481 => "0000011010001011",482 => "0000011010010010",483 => "0000011010011001",
	484 => "0000011010011111",485 => "0000011010100110",486 => "0000011010101100",
	487 => "0000011010110011",488 => "0000011010111010",489 => "0000011011000001",
	490 => "0000011011000111",491 => "0000011011001110",492 => "0000011011010101",
	493 => "0000011011011100",494 => "0000011011100011",495 => "0000011011101010",
	496 => "0000011011110000",497 => "0000011011110111",498 => "0000011011111110",
	499 => "0000011100000101",500 => "0000011100001100",501 => "0000011100010100",
	502 => "0000011100011011",503 => "0000011100100010",504 => "0000011100101001",
	505 => "0000011100110000",506 => "0000011100110111",507 => "0000011100111111",
	508 => "0000011101000110",509 => "0000011101001101",510 => "0000011101010100",
	511 => "0000011101011100",512 => "0000011101100011",513 => "0000011101101011",
	514 => "0000011101110010",515 => "0000011101111001",516 => "0000011110000001",
	517 => "0000011110001000",518 => "0000011110010000",519 => "0000011110011000",
	520 => "0000011110011111",521 => "0000011110100111",522 => "0000011110101110",
	523 => "0000011110110110",524 => "0000011110111110",525 => "0000011111000110",
	526 => "0000011111001101",527 => "0000011111010101",528 => "0000011111011101",
	529 => "0000011111100101",530 => "0000011111101101",531 => "0000011111110101",
	532 => "0000011111111101",533 => "0000100000000101",534 => "0000100000001101",
	535 => "0000100000010101",536 => "0000100000011101",537 => "0000100000100101",
	538 => "0000100000101101",539 => "0000100000110110",540 => "0000100000111110",
	541 => "0000100001000110",542 => "0000100001001110",543 => "0000100001010111",
	544 => "0000100001011111",545 => "0000100001100111",546 => "0000100001110000",
	547 => "0000100001111000",548 => "0000100010000001",549 => "0000100010001001",
	550 => "0000100010010010",551 => "0000100010011010",552 => "0000100010100011",
	553 => "0000100010101100",554 => "0000100010110100",555 => "0000100010111101",
	556 => "0000100011000110",557 => "0000100011001111",558 => "0000100011010111",
	559 => "0000100011100000",560 => "0000100011101001",561 => "0000100011110010",
	562 => "0000100011111011",563 => "0000100100000100",564 => "0000100100001101",
	565 => "0000100100010110",566 => "0000100100011111",567 => "0000100100101000",
	568 => "0000100100110010",569 => "0000100100111011",570 => "0000100101000100",
	571 => "0000100101001101",572 => "0000100101010111",573 => "0000100101100000",
	574 => "0000100101101001",575 => "0000100101110011",576 => "0000100101111100",
	577 => "0000100110000110",578 => "0000100110001111",579 => "0000100110011001",
	580 => "0000100110100011",581 => "0000100110101100",582 => "0000100110110110",
	583 => "0000100111000000",584 => "0000100111001001",585 => "0000100111010011",
	586 => "0000100111011101",587 => "0000100111100111",588 => "0000100111110001",
	589 => "0000100111111011",590 => "0000101000000101",591 => "0000101000001111",
	592 => "0000101000011001",593 => "0000101000100011",594 => "0000101000101101",
	595 => "0000101000110111",596 => "0000101001000010",597 => "0000101001001100",
	598 => "0000101001010110",599 => "0000101001100001",600 => "0000101001101011",
	601 => "0000101001110110",602 => "0000101010000000",603 => "0000101010001011",
	604 => "0000101010010101",605 => "0000101010100000",606 => "0000101010101010",
	607 => "0000101010110101",608 => "0000101011000000",609 => "0000101011001011",
	610 => "0000101011010101",611 => "0000101011100000",612 => "0000101011101011",
	613 => "0000101011110110",614 => "0000101100000001",615 => "0000101100001100",
	616 => "0000101100010111",617 => "0000101100100010",618 => "0000101100101101",
	619 => "0000101100111001",620 => "0000101101000100",621 => "0000101101001111",
	622 => "0000101101011010",623 => "0000101101100110",624 => "0000101101110001",
	625 => "0000101101111101",626 => "0000101110001000",627 => "0000101110010100",
	628 => "0000101110011111",629 => "0000101110101011",630 => "0000101110110111",
	631 => "0000101111000010",632 => "0000101111001110",633 => "0000101111011010",
	634 => "0000101111100110",635 => "0000101111110010",636 => "0000101111111110",
	637 => "0000110000001010",638 => "0000110000010110",639 => "0000110000100010",
	640 => "0000110000101110",641 => "0000110000111010",642 => "0000110001000111",
	643 => "0000110001010011",644 => "0000110001011111",645 => "0000110001101100",
	646 => "0000110001111000",647 => "0000110010000101",648 => "0000110010010001",
	649 => "0000110010011110",650 => "0000110010101010",651 => "0000110010110111",
	652 => "0000110011000100",653 => "0000110011010001",654 => "0000110011011110",
	655 => "0000110011101010",656 => "0000110011110111",657 => "0000110100000100",
	658 => "0000110100010001",659 => "0000110100011110",660 => "0000110100101100",
	661 => "0000110100111001",662 => "0000110101000110",663 => "0000110101010011",
	664 => "0000110101100001",665 => "0000110101101110",666 => "0000110101111100",
	667 => "0000110110001001",668 => "0000110110010111",669 => "0000110110100100",
	670 => "0000110110110010",671 => "0000110111000000",672 => "0000110111001101",
	673 => "0000110111011011",674 => "0000110111101001",675 => "0000110111110111",
	676 => "0000111000000101",677 => "0000111000010011",678 => "0000111000100001",
	679 => "0000111000101111",680 => "0000111000111110",681 => "0000111001001100",
	682 => "0000111001011010",683 => "0000111001101001",684 => "0000111001110111",
	685 => "0000111010000110",686 => "0000111010010100",687 => "0000111010100011",
	688 => "0000111010110001",689 => "0000111011000000",690 => "0000111011001111",
	691 => "0000111011011110",692 => "0000111011101101",693 => "0000111011111100",
	694 => "0000111100001011",695 => "0000111100011010",696 => "0000111100101001",
	697 => "0000111100111000",698 => "0000111101000111",699 => "0000111101010111",
	700 => "0000111101100110",701 => "0000111101110101",702 => "0000111110000101",
	703 => "0000111110010100",704 => "0000111110100100",705 => "0000111110110100",
	706 => "0000111111000011",707 => "0000111111010011",708 => "0000111111100011",
	709 => "0000111111110011",710 => "0001000000000011",711 => "0001000000010011",
	712 => "0001000000100011",713 => "0001000000110011",714 => "0001000001000100",
	715 => "0001000001010100",716 => "0001000001100100",717 => "0001000001110101",
	718 => "0001000010000101",719 => "0001000010010110",720 => "0001000010100110",
	721 => "0001000010110111",722 => "0001000011001000",723 => "0001000011011001",
	724 => "0001000011101001",725 => "0001000011111010",726 => "0001000100001011",
	727 => "0001000100011100",728 => "0001000100101110",729 => "0001000100111111",
	730 => "0001000101010000",731 => "0001000101100001",732 => "0001000101110011",
	733 => "0001000110000100",734 => "0001000110010110",735 => "0001000110101000",
	736 => "0001000110111001",737 => "0001000111001011",738 => "0001000111011101",
	739 => "0001000111101111",740 => "0001001000000001",741 => "0001001000010011",
	742 => "0001001000100101",743 => "0001001000110111",744 => "0001001001001001",
	745 => "0001001001011100",746 => "0001001001101110",747 => "0001001010000000",
	748 => "0001001010010011",749 => "0001001010100110",750 => "0001001010111000",
	751 => "0001001011001011",752 => "0001001011011110",753 => "0001001011110001",
	754 => "0001001100000100",755 => "0001001100010111",756 => "0001001100101010",
	757 => "0001001100111101",758 => "0001001101010000",759 => "0001001101100100",
	760 => "0001001101110111",761 => "0001001110001011",762 => "0001001110011110",
	763 => "0001001110110010",764 => "0001001111000110",765 => "0001001111011001",
	766 => "0001001111101101",767 => "0001010000000001",768 => "0001010000010101",
	769 => "0001010000101010",770 => "0001010000111110",771 => "0001010001010010",
	772 => "0001010001100110",773 => "0001010001111011",774 => "0001010010001111",
	775 => "0001010010100100",776 => "0001010010111001",777 => "0001010011001101",
	778 => "0001010011100010",779 => "0001010011110111",780 => "0001010100001100",
	781 => "0001010100100001",782 => "0001010100110110",783 => "0001010101001100",
	784 => "0001010101100001",785 => "0001010101110110",786 => "0001010110001100",
	787 => "0001010110100010",788 => "0001010110110111",789 => "0001010111001101",
	790 => "0001010111100011",791 => "0001010111111001",792 => "0001011000001111",
	793 => "0001011000100101",794 => "0001011000111011",795 => "0001011001010001",
	796 => "0001011001101000",797 => "0001011001111110",798 => "0001011010010101",
	799 => "0001011010101011",800 => "0001011011000010",801 => "0001011011011001",
	802 => "0001011011110000",803 => "0001011100000111",804 => "0001011100011110",
	805 => "0001011100110101",806 => "0001011101001100",807 => "0001011101100100",
	808 => "0001011101111011",809 => "0001011110010011",810 => "0001011110101010",
	811 => "0001011111000010",812 => "0001011111011010",813 => "0001011111110010",
	814 => "0001100000001010",815 => "0001100000100010",816 => "0001100000111010",
	817 => "0001100001010010",818 => "0001100001101010",819 => "0001100010000011",
	820 => "0001100010011011",821 => "0001100010110100",822 => "0001100011001101",
	823 => "0001100011100110",824 => "0001100011111111",825 => "0001100100011000",
	826 => "0001100100110001",827 => "0001100101001010",828 => "0001100101100011",
	829 => "0001100101111101",830 => "0001100110010110",831 => "0001100110110000",
	832 => "0001100111001010",833 => "0001100111100100",834 => "0001100111111110",
	835 => "0001101000011000",836 => "0001101000110010",837 => "0001101001001100",
	838 => "0001101001100110",839 => "0001101010000001",840 => "0001101010011011",
	841 => "0001101010110110",842 => "0001101011010001",843 => "0001101011101100",
	844 => "0001101100000111",845 => "0001101100100010",846 => "0001101100111101",
	847 => "0001101101011000",848 => "0001101101110100",849 => "0001101110001111",
	850 => "0001101110101011",851 => "0001101111000110",852 => "0001101111100010",
	853 => "0001101111111110",854 => "0001110000011010",855 => "0001110000110110",
	856 => "0001110001010011",857 => "0001110001101111",858 => "0001110010001100",
	859 => "0001110010101000",860 => "0001110011000101",861 => "0001110011100010",
	862 => "0001110011111111",863 => "0001110100011100",864 => "0001110100111001",
	865 => "0001110101010110",866 => "0001110101110100",867 => "0001110110010001",
	868 => "0001110110101111",869 => "0001110111001100",870 => "0001110111101010",
	871 => "0001111000001000",872 => "0001111000100110",873 => "0001111001000101",
	874 => "0001111001100011",875 => "0001111010000001",876 => "0001111010100000",
	877 => "0001111010111111",878 => "0001111011011101",879 => "0001111011111100",
	880 => "0001111100011011",881 => "0001111100111011",882 => "0001111101011010",
	883 => "0001111101111001",884 => "0001111110011001",885 => "0001111110111001",
	886 => "0001111111011000",887 => "0001111111111000",888 => "0010000000011000",
	889 => "0010000000111000",890 => "0010000001011001",891 => "0010000001111001",
	892 => "0010000010011010",893 => "0010000010111010",894 => "0010000011011011",
	895 => "0010000011111100",896 => "0010000100011101",897 => "0010000100111110",
	898 => "0010000101100000",899 => "0010000110000001",900 => "0010000110100011",
	901 => "0010000111000100",902 => "0010000111100110",903 => "0010001000001000",
	904 => "0010001000101010",905 => "0010001001001100",906 => "0010001001101111",
	907 => "0010001010010001",908 => "0010001010110100",909 => "0010001011010111",
	910 => "0010001011111010",911 => "0010001100011101",912 => "0010001101000000",
	913 => "0010001101100011",914 => "0010001110000111",915 => "0010001110101010",
	916 => "0010001111001110",917 => "0010001111110010",918 => "0010010000010110",
	919 => "0010010000111010",920 => "0010010001011110",921 => "0010010010000011",
	922 => "0010010010100111",923 => "0010010011001100",924 => "0010010011110001",
	925 => "0010010100010110",926 => "0010010100111011",927 => "0010010101100000",
	928 => "0010010110000110",929 => "0010010110101011",930 => "0010010111010001",
	931 => "0010010111110111",932 => "0010011000011101",933 => "0010011001000011",
	934 => "0010011001101010",935 => "0010011010010000",936 => "0010011010110111",
	937 => "0010011011011110",938 => "0010011100000101",939 => "0010011100101100",
	940 => "0010011101010011",941 => "0010011101111010",942 => "0010011110100010",
	943 => "0010011111001010",944 => "0010011111110001",945 => "0010100000011001",
	946 => "0010100001000010",947 => "0010100001101010",948 => "0010100010010010",
	949 => "0010100010111011",950 => "0010100011100100",951 => "0010100100001101",
	952 => "0010100100110110",953 => "0010100101011111",954 => "0010100110001001",
	955 => "0010100110110010",956 => "0010100111011100",957 => "0010101000000110",
	958 => "0010101000110000",959 => "0010101001011010",960 => "0010101010000101",
	961 => "0010101010110000",962 => "0010101011011010",963 => "0010101100000101",
	964 => "0010101100110000",965 => "0010101101011100",966 => "0010101110000111",
	967 => "0010101110110011",968 => "0010101111011110",969 => "0010110000001010",
	970 => "0010110000110111",971 => "0010110001100011",972 => "0010110010001111",
	973 => "0010110010111100",974 => "0010110011101001",975 => "0010110100010110",
	976 => "0010110101000011",977 => "0010110101110000",978 => "0010110110011110",
	979 => "0010110111001100",980 => "0010110111111001",981 => "0010111000100111",
	982 => "0010111001010110",983 => "0010111010000100",984 => "0010111010110011",
	985 => "0010111011100010",986 => "0010111100010001",987 => "0010111101000000",
	988 => "0010111101101111",989 => "0010111110011111",990 => "0010111111001110",
	991 => "0010111111111110",992 => "0011000000101110",993 => "0011000001011111",
	994 => "0011000010001111",995 => "0011000011000000",996 => "0011000011110001",
	997 => "0011000100100010",998 => "0011000101010011",999 => "0011000110000100",
	1000 => "0011000110110110",1001 => "0011000111101000",1002 => "0011001000011010",
	1003 => "0011001001001100",1004 => "0011001001111110",1005 => "0011001010110001",
	1006 => "0011001011100100",1007 => "0011001100010111",1008 => "0011001101001010",
	1009 => "0011001101111101",1010 => "0011001110110001",1011 => "0011001111100101",
	1012 => "0011010000011001",1013 => "0011010001001101",1014 => "0011010010000001",
	1015 => "0011010010110110",1016 => "0011010011101011",1017 => "0011010100100000",
	1018 => "0011010101010101",1019 => "0011010110001010",1020 => "0011010111000000",
	1021 => "0011010111110110",1022 => "0011011000101100",1023 => "0011011001100010",
	1024 => "0011011010011001",1025 => "0011011011001111",1026 => "0011011100000110",
	1027 => "0011011100111101",1028 => "0011011101110101",1029 => "0011011110101100",
	1030 => "0011011111100100",1031 => "0011100000011100",1032 => "0011100001010100",
	1033 => "0011100010001101",1034 => "0011100011000101",1035 => "0011100011111110",
	1036 => "0011100100110111",1037 => "0011100101110001",1038 => "0011100110101010",
	1039 => "0011100111100100",1040 => "0011101000011110",1041 => "0011101001011000",
	1042 => "0011101010010011",1043 => "0011101011001101",1044 => "0011101100001000",
	1045 => "0011101101000100",1046 => "0011101101111111",1047 => "0011101110111011",
	1048 => "0011101111110110",1049 => "0011110000110010",1050 => "0011110001101111",
	1051 => "0011110010101011",1052 => "0011110011101000",1053 => "0011110100100101",
	1054 => "0011110101100010",1055 => "0011110110100000",1056 => "0011110111011110",
	1057 => "0011111000011100",1058 => "0011111001011010",1059 => "0011111010011000",
	1060 => "0011111011010111",1061 => "0011111100010110",1062 => "0011111101010101",
	1063 => "0011111110010101",1064 => "0011111111010100",1065 => "0100000000010100",
	1066 => "0100000001010101",1067 => "0100000010010101",1068 => "0100000011010110",
	1069 => "0100000100010111",1070 => "0100000101011000",1071 => "0100000110011001",
	1072 => "0100000111011011",1073 => "0100001000011101",1074 => "0100001001011111",
	1075 => "0100001010100010",1076 => "0100001011100101",1077 => "0100001100101000",
	1078 => "0100001101101011",1079 => "0100001110101110",1080 => "0100001111110010",
	1081 => "0100010000110110",1082 => "0100010001111011",1083 => "0100010010111111",
	1084 => "0100010100000100",1085 => "0100010101001001",1086 => "0100010110001111",
	1087 => "0100010111010101",1088 => "0100011000011010",1089 => "0100011001100001",
	1090 => "0100011010100111",1091 => "0100011011101110",1092 => "0100011100110101",
	1093 => "0100011101111100",1094 => "0100011111000100",1095 => "0100100000001100",
	1096 => "0100100001010100",1097 => "0100100010011101",1098 => "0100100011100101",
	1099 => "0100100100101110",1100 => "0100100101111000",1101 => "0100100111000001",
	1102 => "0100101000001011",1103 => "0100101001010101",1104 => "0100101010100000",
	1105 => "0100101011101011",1106 => "0100101100110110",1107 => "0100101110000001",
	1108 => "0100101111001101",1109 => "0100110000011001",1110 => "0100110001100101",
	1111 => "0100110010110010",1112 => "0100110011111110",1113 => "0100110101001100",
	1114 => "0100110110011001",1115 => "0100110111100111",1116 => "0100111000110101",
	1117 => "0100111010000011",1118 => "0100111011010010",1119 => "0100111100100001",
	1120 => "0100111101110000",1121 => "0100111111000000",1122 => "0101000000010000",
	1123 => "0101000001100000",1124 => "0101000010110000",1125 => "0101000100000001",
	1126 => "0101000101010010",1127 => "0101000110100100",1128 => "0101000111110110",
	1129 => "0101001001001000",1130 => "0101001010011010",1131 => "0101001011101101",
	1132 => "0101001101000000",1133 => "0101001110010011",1134 => "0101001111100111",
	1135 => "0101010000111011",1136 => "0101010010010000",1137 => "0101010011100100",
	1138 => "0101010100111001",1139 => "0101010110001111",1140 => "0101010111100101",
	1141 => "0101011000111011",1142 => "0101011010010001",1143 => "0101011011101000",
	1144 => "0101011100111111",1145 => "0101011110010110",1146 => "0101011111101110",
	1147 => "0101100001000110",1148 => "0101100010011111",1149 => "0101100011110111",
	1150 => "0101100101010001",1151 => "0101100110101010",1152 => "0101101000000100",
	1153 => "0101101001011110",1154 => "0101101010111001",1155 => "0101101100010100",
	1156 => "0101101101101111",1157 => "0101101111001010",1158 => "0101110000100110",
	1159 => "0101110010000011",1160 => "0101110011011111",1161 => "0101110100111100",
	1162 => "0101110110011010",1163 => "0101110111111000",1164 => "0101111001010110",
	1165 => "0101111010110100",1166 => "0101111100010011",1167 => "0101111101110010",
	1168 => "0101111111010010",1169 => "0110000000110010",1170 => "0110000010010011",
	1171 => "0110000011110011",1172 => "0110000101010100",1173 => "0110000110110110",
	1174 => "0110001000011000",1175 => "0110001001111010",1176 => "0110001011011101",
	1177 => "0110001101000000",1178 => "0110001110100011",1179 => "0110010000000111",
	1180 => "0110010001101011",1181 => "0110010011010000",1182 => "0110010100110101",
	1183 => "0110010110011010",1184 => "0110011000000000",1185 => "0110011001100110",
	1186 => "0110011011001101",1187 => "0110011100110100",1188 => "0110011110011011",
	1189 => "0110100000000011",1190 => "0110100001101011",1191 => "0110100011010100",
	1192 => "0110100100111101",1193 => "0110100110100111",1194 => "0110101000010000",
	1195 => "0110101001111011",1196 => "0110101011100101",1197 => "0110101101010000",
	1198 => "0110101110111100",1199 => "0110110000101000",1200 => "0110110010010100",
	1201 => "0110110100000001",1202 => "0110110101101110",1203 => "0110110111011100",
	1204 => "0110111001001010",1205 => "0110111010111001",1206 => "0110111100101000",
	1207 => "0110111110010111",1208 => "0111000000000111",1209 => "0111000001110111",
	1210 => "0111000011101000",1211 => "0111000101011001",1212 => "0111000111001010",
	1213 => "0111001000111100",1214 => "0111001010101111",1215 => "0111001100100010",
	1216 => "0111001110010101",1217 => "0111010000001001",1218 => "0111010001111101",
	1219 => "0111010011110010",1220 => "0111010101100111",1221 => "0111010111011101",
	1222 => "0111011001010011",1223 => "0111011011001001",1224 => "0111011101000000",
	1225 => "0111011110111000",1226 => "0111100000110000",1227 => "0111100010101000",
	1228 => "0111100100100001",1229 => "0111100110011010",1230 => "0111101000010100",
	1231 => "0111101010001111",1232 => "0111101100001001",1233 => "0111101110000101",
	1234 => "0111110000000000",1235 => "0111110001111101",1236 => "0111110011111001",
	1237 => "0111110101110111",1238 => "0111110111110100",1239 => "0111111001110011",
	1240 => "0111111011110001",1241 => "0111111101110000",1242 => "0000000000000000",
	1243 => "0000000000000000",1244 => "0000000000000000",1245 => "0000000000000000",
	1246 => "0000000000000000",1247 => "0000000000000000",1248 => "0000000000000000",
	1249 => "0000000000000000",1250 => "0000000000000000",1251 => "0000000000000000",
	1252 => "0000000000000000",1253 => "0000000000000000",1254 => "0000000000000000",
	1255 => "0000000000000000",1256 => "0000000000000000",1257 => "0000000000000000",
	1258 => "0000000000000000",1259 => "0000000000000000",1260 => "0000000000000000",
	1261 => "0000000000000000",1262 => "0000000000000000",1263 => "0000000000000000",
	1264 => "0000000000000000",1265 => "0000000000000000",1266 => "0000000000000000",
	1267 => "0000000000000000",1268 => "0000000000000000",1269 => "0000000000000000",
	1270 => "0000000000000000",1271 => "0000000000000000",1272 => "0000000000000000",
	1273 => "0000000000000000",1274 => "0000000000000000",1275 => "0000000000000000",
	1276 => "0000000000000000",1277 => "0000000000000000",1278 => "0000000000000000",
	1279 => "0000000000000000",1280 => "0000000000000000",1281 => "0000000000000000",
	1282 => "0000000000000000",1283 => "0000000000000000",1284 => "0000000000000000",
	1285 => "0000000000000000",1286 => "0000000000000000",1287 => "0000000000000000",
	1288 => "0000000000000000",1289 => "0000000000000000",1290 => "0000000000000000",
	1291 => "0000000000000000",1292 => "0000000000000000",1293 => "0000000000000000",
	1294 => "0000000000000000",1295 => "0000000000000000",1296 => "0000000000000000",
	1297 => "0000000000000000",1298 => "0000000000000000",1299 => "0000000000000000",
	1300 => "0000000000000000",1301 => "0000000000000000",1302 => "0000000000000000",
	1303 => "0000000000000000",1304 => "0000000000000000",1305 => "0000000000000000",
	1306 => "0000000000000000",1307 => "0000000000000000",1308 => "0000000000000000",
	1309 => "0000000000000000",1310 => "0000000000000000",1311 => "0000000000000000",
	1312 => "0000000000000000",1313 => "0000000000000000",1314 => "0000000000000000",
	1315 => "0000000000000000",1316 => "0000000000000000",1317 => "0000000000000000",
	1318 => "0000000000000000",1319 => "0000000000000000",1320 => "0000000000000000",
	1321 => "0000000000000000",1322 => "0000000000000000",1323 => "0000000000000000",
	1324 => "0000000000000000",1325 => "0000000000000000",1326 => "0000000000000000",
	1327 => "0000000000000000",1328 => "0000000000000000",1329 => "0000000000000000",
	1330 => "0000000000000000",1331 => "0000000000000000",1332 => "0000000000000000",
	1333 => "0000000000000000",1334 => "0000000000000000",1335 => "0000000000000000",
	1336 => "0000000000000000",1337 => "0000000000000000",1338 => "0000000000000000",
	1339 => "0000000000000000",1340 => "0000000000000000",1341 => "0000000000000000",
	1342 => "0000000000000000",1343 => "0000000000000000",1344 => "0000000000000000",
	1345 => "0000000000000000",1346 => "0000000000000000",1347 => "0000000000000000",
	1348 => "0000000000000000",1349 => "0000000000000000",1350 => "0000000000000000",
	1351 => "0000000000000000",1352 => "0000000000000000",1353 => "0000000000000000",
	1354 => "0000000000000000",1355 => "0000000000000000",1356 => "0000000000000000",
	1357 => "0000000000000000",1358 => "0000000000000000",1359 => "0000000000000000",
	1360 => "0000000000000000",1361 => "0000000000000000",1362 => "0000000000000000",
	1363 => "0000000000000000",1364 => "0000000000000000",1365 => "0000000000000000",
	1366 => "0000000000000000",1367 => "0000000000000000",1368 => "0000000000000000",
	1369 => "0000000000000000",1370 => "0000000000000000",1371 => "0000000000000000",
	1372 => "0000000000000000",1373 => "0000000000000000",1374 => "0000000000000000",
	1375 => "0000000000000000",1376 => "0000000000000000",1377 => "0000000000000000",
	1378 => "0000000000000000",1379 => "0000000000000000",1380 => "0000000000000000",
	1381 => "0000000000000000",1382 => "0000000000000000",1383 => "0000000000000000",
	1384 => "0000000000000000",1385 => "0000000000000000",1386 => "0000000000000000",
	1387 => "0000000000000000",1388 => "0000000000000000",1389 => "0000000000000000",
	1390 => "0000000000000000",1391 => "0000000000000000",1392 => "0000000000000000",
	1393 => "0000000000000000",1394 => "0000000000000000",1395 => "0000000000000000",
	1396 => "0000000000000000",1397 => "0000000000000000",1398 => "0000000000000000",
	1399 => "0000000000000000",1400 => "0000000000000000",1401 => "0000000000000000",
	1402 => "0000000000000000",1403 => "0000000000000000",1404 => "0000000000000000",
	1405 => "0000000000000000",1406 => "0000000000000000",1407 => "0000000000000000",
	1408 => "0000000000000000",1409 => "0000000000000000",1410 => "0000000000000000",
	1411 => "0000000000000000",1412 => "0000000000000000",1413 => "0000000000000000",
	1414 => "0000000000000000",1415 => "0000000000000000",1416 => "0000000000000000",
	1417 => "0000000000000000",1418 => "0000000000000000",1419 => "0000000000000000",
	1420 => "0000000000000000",1421 => "0000000000000000",1422 => "0000000000000000",
	1423 => "0000000000000000",1424 => "0000000000000000",1425 => "0000000000000000",
	1426 => "0000000000000000",1427 => "0000000000000000",1428 => "0000000000000000",
	1429 => "0000000000000000",1430 => "0000000000000000",1431 => "0000000000000000",
	1432 => "0000000000000000",1433 => "0000000000000000",1434 => "0000000000000000",
	1435 => "0000000000000000",1436 => "0000000000000000",1437 => "0000000000000000",
	1438 => "0000000000000000",1439 => "0000000000000000",1440 => "0000000000000000",
	1441 => "0000000000000000",1442 => "0000000000000000",1443 => "0000000000000000",
	1444 => "0000000000000000",1445 => "0000000000000000",1446 => "0000000000000000",
	1447 => "0000000000000000",1448 => "0000000000000000",1449 => "0000000000000000",
	1450 => "0000000000000000",1451 => "0000000000000000",1452 => "0000000000000000",
	1453 => "0000000000000000",1454 => "0000000000000000",1455 => "0000000000000000",
	1456 => "0000000000000000",1457 => "0000000000000000",1458 => "0000000000000000",
	1459 => "0000000000000000",1460 => "0000000000000000",1461 => "0000000000000000",
	1462 => "0000000000000000",1463 => "0000000000000000",1464 => "0000000000000000",
	1465 => "0000000000000000",1466 => "0000000000000000",1467 => "0000000000000000",
	1468 => "0000000000000000",1469 => "0000000000000000",1470 => "0000000000000000",
	1471 => "0000000000000000",1472 => "0000000000000000",1473 => "0000000000000000",
	1474 => "0000000000000000",1475 => "0000000000000000",1476 => "0000000000000000",
	1477 => "0000000000000000",1478 => "0000000000000000",1479 => "0000000000000000",
	1480 => "0000000000000000",1481 => "0000000000000000",1482 => "0000000000000000",
	1483 => "0000000000000000",1484 => "0000000000000000",1485 => "0000000000000000",
	1486 => "0000000000000000",1487 => "0000000000000000",1488 => "0000000000000000",
	1489 => "0000000000000000",1490 => "0000000000000000",1491 => "0000000000000000",
	1492 => "0000000000000000",1493 => "0000000000000000",1494 => "0000000000000000",
	1495 => "0000000000000000",1496 => "0000000000000000",1497 => "0000000000000000",
	1498 => "0000000000000000",1499 => "0000000000000000",1500 => "0000000000000000",
	1501 => "0000000000000000",1502 => "0000000000000000",1503 => "0000000000000000",
	1504 => "0000000000000000",1505 => "0000000000000000",1506 => "0000000000000000",
	1507 => "0000000000000000",1508 => "0000000000000000",1509 => "0000000000000000",
	1510 => "0000000000000000",1511 => "0000000000000000",1512 => "0000000000000000",
	1513 => "0000000000000000",1514 => "0000000000000000",1515 => "0000000000000000",
	1516 => "0000000000000000",1517 => "0000000000000000",1518 => "0000000000000000",
	1519 => "0000000000000000",1520 => "0000000000000000",1521 => "0000000000000000",
	1522 => "0000000000000000",1523 => "0000000000000000",1524 => "0000000000000000",
	1525 => "0000000000000000",1526 => "0000000000000000",1527 => "0000000000000000",
	1528 => "0000000000000000",1529 => "0000000000000000",1530 => "0000000000000000",
	1531 => "0000000000000000",1532 => "0000000000000000",1533 => "0000000000000000",
	1534 => "0000000000000000",1535 => "0000000000000000",1536 => "0000000000000000",
	1537 => "0000000000000000",1538 => "0000000000000000",1539 => "0000000000000000",
	1540 => "0000000000000000",1541 => "0000000000000000",1542 => "0000000000000000",
	1543 => "0000000000000000",1544 => "0000000000000000",1545 => "0000000000000000",
	1546 => "0000000000000000",1547 => "0000000000000000",1548 => "0000000000000000",
	1549 => "0000000000000000",1550 => "0000000000000000",1551 => "0000000000000000",
	1552 => "0000000000000000",1553 => "0000000000000000",1554 => "0000000000000000",
	1555 => "0000000000000000",1556 => "0000000000000000",1557 => "0000000000000000",
	1558 => "0000000000000000",1559 => "0000000000000000",1560 => "0000000000000000",
	1561 => "0000000000000000",1562 => "0000000000000000",1563 => "0000000000000000",
	1564 => "0000000000000000",1565 => "0000000000000000",1566 => "0000000000000000",
	1567 => "0000000000000000",1568 => "0000000000000000",1569 => "0000000000000000",
	1570 => "0000000000000000",1571 => "0000000000000000",1572 => "0000000000000000",
	1573 => "0000000000000000",1574 => "0000000000000000",1575 => "0000000000000000",
	1576 => "0000000000000000",1577 => "0000000000000000",1578 => "0000000000000000",
	1579 => "0000000000000000",1580 => "0000000000000000",1581 => "0000000000000000",
	1582 => "0000000000000000",1583 => "0000000000000000",1584 => "0000000000000000",
	1585 => "0000000000000000",1586 => "0000000000000000",1587 => "0000000000000000",
	1588 => "0000000000000000",1589 => "0000000000000000",1590 => "0000000000000000",
	1591 => "0000000000000000",1592 => "0000000000000000",1593 => "0000000000000000",
	1594 => "0000000000000000",1595 => "0000000000000000",1596 => "0000000000000000",
	1597 => "0000000000000000",1598 => "0000000000000000",1599 => "0000000000000000",
	1600 => "0000000000000000",1601 => "0000000000000000",1602 => "0000000000000000",
	1603 => "0000000000000000",1604 => "0000000000000000",1605 => "0000000000000000",
	1606 => "0000000000000000",1607 => "0000000000000000",1608 => "0000000000000000",
	1609 => "0000000000000000",1610 => "0000000000000000",1611 => "0000000000000000",
	1612 => "0000000000000000",1613 => "0000000000000000",1614 => "0000000000000000",
	1615 => "0000000000000000",1616 => "0000000000000000",1617 => "0000000000000000",
	1618 => "0000000000000000",1619 => "0000000000000000",1620 => "0000000000000000",
	1621 => "0000000000000000",1622 => "0000000000000000",1623 => "0000000000000000",
	1624 => "0000000000000000",1625 => "0000000000000000",1626 => "0000000000000000",
	1627 => "0000000000000000",1628 => "0000000000000000",1629 => "0000000000000000",
	1630 => "0000000000000000",1631 => "0000000000000000",1632 => "0000000000000000",
	1633 => "0000000000000000",1634 => "0000000000000000",1635 => "0000000000000000",
	1636 => "0000000000000000",1637 => "0000000000000000",1638 => "0000000000000000",
	1639 => "0000000000000000",1640 => "0000000000000000",1641 => "0000000000000000",
	1642 => "0000000000000000",1643 => "0000000000000000",1644 => "0000000000000000",
	1645 => "0000000000000000",1646 => "0000000000000000",1647 => "0000000000000000",
	1648 => "0000000000000000",1649 => "0000000000000000",1650 => "0000000000000000",
	1651 => "0000000000000000",1652 => "0000000000000000",1653 => "0000000000000000",
	1654 => "0000000000000000",1655 => "0000000000000000",1656 => "0000000000000000",
	1657 => "0000000000000000",1658 => "0000000000000000",1659 => "0000000000000000",
	1660 => "0000000000000000",1661 => "0000000000000000",1662 => "0000000000000000",
	1663 => "0000000000000000",1664 => "0000000000000000",1665 => "0000000000000000",
	1666 => "0000000000000000",1667 => "0000000000000000",1668 => "0000000000000000",
	1669 => "0000000000000000",1670 => "0000000000000000",1671 => "0000000000000000",
	1672 => "0000000000000000",1673 => "0000000000000000",1674 => "0000000000000000",
	1675 => "0000000000000000",1676 => "0000000000000000",1677 => "0000000000000000",
	1678 => "0000000000000000",1679 => "0000000000000000",1680 => "0000000000000000",
	1681 => "0000000000000000",1682 => "0000000000000000",1683 => "0000000000000000",
	1684 => "0000000000000000",1685 => "0000000000000000",1686 => "0000000000000000",
	1687 => "0000000000000000",1688 => "0000000000000000",1689 => "0000000000000000",
	1690 => "0000000000000000",1691 => "0000000000000000",1692 => "0000000000000000",
	1693 => "0000000000000000",1694 => "0000000000000000",1695 => "0000000000000000",
	1696 => "0000000000000000",1697 => "0000000000000000",1698 => "0000000000000000",
	1699 => "0000000000000000",1700 => "0000000000000000",1701 => "0000000000000000",
	1702 => "0000000000000000",1703 => "0000000000000000",1704 => "0000000000000000",
	1705 => "0000000000000000",1706 => "0000000000000000",1707 => "0000000000000000",
	1708 => "0000000000000000",1709 => "0000000000000000",1710 => "0000000000000000",
	1711 => "0000000000000000",1712 => "0000000000000000",1713 => "0000000000000000",
	1714 => "0000000000000000",1715 => "0000000000000000",1716 => "0000000000000000",
	1717 => "0000000000000000",1718 => "0000000000000000",1719 => "0000000000000000",
	1720 => "0000000000000000",1721 => "0000000000000000",1722 => "0000000000000000",
	1723 => "0000000000000000",1724 => "0000000000000000",1725 => "0000000000000000",
	1726 => "0000000000000000",1727 => "0000000000000000",1728 => "0000000000000000",
	1729 => "0000000000000000",1730 => "0000000000000000",1731 => "0000000000000000",
	1732 => "0000000000000000",1733 => "0000000000000000",1734 => "0000000000000000",
	1735 => "0000000000000000",1736 => "0000000000000000",1737 => "0000000000000000",
	1738 => "0000000000000000",1739 => "0000000000000000",1740 => "0000000000000000",
	1741 => "0000000000000000",1742 => "0000000000000000",1743 => "0000000000000000",
	1744 => "0000000000000000",1745 => "0000000000000000",1746 => "0000000000000000",
	1747 => "0000000000000000",1748 => "0000000000000000",1749 => "0000000000000000",
	1750 => "0000000000000000",1751 => "0000000000000000",1752 => "0000000000000000",
	1753 => "0000000000000000",1754 => "0000000000000000",1755 => "0000000000000000",
	1756 => "0000000000000000",1757 => "0000000000000000",1758 => "0000000000000000",
	1759 => "0000000000000000",1760 => "0000000000000000",1761 => "0000000000000000",
	1762 => "0000000000000000",1763 => "0000000000000000",1764 => "0000000000000000",
	1765 => "0000000000000000",1766 => "0000000000000000",1767 => "0000000000000000",
	1768 => "0000000000000000",1769 => "0000000000000000",1770 => "0000000000000000",
	1771 => "0000000000000000",1772 => "0000000000000000",1773 => "0000000000000000",
	1774 => "0000000000000000",1775 => "0000000000000000",1776 => "0000000000000000",
	1777 => "0000000000000000",1778 => "0000000000000000",1779 => "0000000000000000",
	1780 => "0000000000000000",1781 => "0000000000000000",1782 => "0000000000000000",
	1783 => "0000000000000000",1784 => "0000000000000000",1785 => "0000000000000000",
	1786 => "0000000000000000",1787 => "0000000000000000",1788 => "0000000000000000",
	1789 => "0000000000000000",1790 => "0000000000000000",1791 => "0000000000000000",
	1792 => "0000000000000000",1793 => "0000000000000000",1794 => "0000000000000000",
	1795 => "0000000000000000",1796 => "0000000000000000",1797 => "0000000000000000",
	1798 => "0000000000000000",1799 => "0000000000000000",1800 => "0000000000000000",
	1801 => "0000000000000000",1802 => "0000000000000000",1803 => "0000000000000000",
	1804 => "0000000000000000",1805 => "0000000000000000",1806 => "0000000000000000",
	1807 => "0000000000000000",1808 => "0000000000000000",1809 => "0000000000000000",
	1810 => "0000000000000000",1811 => "0000000000000000",1812 => "0000000000000000",
	1813 => "0000000000000000",1814 => "0000000000000000",1815 => "0000000000000000",
	1816 => "0000000000000000",1817 => "0000000000000000",1818 => "0000000000000000",
	1819 => "0000000000000000",1820 => "0000000000000000",1821 => "0000000000000000",
	1822 => "0000000000000000",1823 => "0000000000000000",1824 => "0000000000000000",
	1825 => "0000000000000000",1826 => "0000000000000000",1827 => "0000000000000000",
	1828 => "0000000000000000",1829 => "0000000000000000",1830 => "0000000000000000",
	1831 => "0000000000000000",1832 => "0000000000000000",1833 => "0000000000000000",
	1834 => "0000000000000000",1835 => "0000000000000000",1836 => "0000000000000000",
	1837 => "0000000000000000",1838 => "0000000000000000",1839 => "0000000000000000",
	1840 => "0000000000000000",1841 => "0000000000000000",1842 => "0000000000000000",
	1843 => "0000000000000000",1844 => "0000000000000000",1845 => "0000000000000000",
	1846 => "0000000000000000",1847 => "0000000000000000",1848 => "0000000000000000",
	1849 => "0000000000000000",1850 => "0000000000000000",1851 => "0000000000000000",
	1852 => "0000000000000000",1853 => "0000000000000000",1854 => "0000000000000000",
	1855 => "0000000000000000",1856 => "0000000000000000",1857 => "0000000000000000",
	1858 => "0000000000000000",1859 => "0000000000000000",1860 => "0000000000000000",
	1861 => "0000000000000000",1862 => "0000000000000000",1863 => "0000000000000000",
	1864 => "0000000000000000",1865 => "0000000000000000",1866 => "0000000000000000",
	1867 => "0000000000000000",1868 => "0000000000000000",1869 => "0000000000000000",
	1870 => "0000000000000000",1871 => "0000000000000000",1872 => "0000000000000000",
	1873 => "0000000000000000",1874 => "0000000000000000",1875 => "0000000000000000",
	1876 => "0000000000000000",1877 => "0000000000000000",1878 => "0000000000000000",
	1879 => "0000000000000000",1880 => "0000000000000000",1881 => "0000000000000000",
	1882 => "0000000000000000",1883 => "0000000000000000",1884 => "0000000000000000",
	1885 => "0000000000000000",1886 => "0000000000000000",1887 => "0000000000000000",
	1888 => "0000000000000000",1889 => "0000000000000000",1890 => "0000000000000000",
	1891 => "0000000000000000",1892 => "0000000000000000",1893 => "0000000000000000",
	1894 => "0000000000000000",1895 => "0000000000000000",1896 => "0000000000000000",
	1897 => "0000000000000000",1898 => "0000000000000000",1899 => "0000000000000000",
	1900 => "0000000000000000",1901 => "0000000000000000",1902 => "0000000000000000",
	1903 => "0000000000000000",1904 => "0000000000000000",1905 => "0000000000000000",
	1906 => "0000000000000000",1907 => "0000000000000000",1908 => "0000000000000000",
	1909 => "0000000000000000",1910 => "0000000000000000",1911 => "0000000000000000",
	1912 => "0000000000000000",1913 => "0000000000000000",1914 => "0000000000000000",
	1915 => "0000000000000000",1916 => "0000000000000000",1917 => "0000000000000000",
	1918 => "0000000000000000",1919 => "0000000000000000",1920 => "0000000000000000",
	1921 => "0000000000000000",1922 => "0000000000000000",1923 => "0000000000000000",
	1924 => "0000000000000000",1925 => "0000000000000000",1926 => "0000000000000000",
	1927 => "0000000000000000",1928 => "0000000000000000",1929 => "0000000000000000",
	1930 => "0000000000000000",1931 => "0000000000000000",1932 => "0000000000000000",
	1933 => "0000000000000000",1934 => "0000000000000000",1935 => "0000000000000000",
	1936 => "0000000000000000",1937 => "0000000000000000",1938 => "0000000000000000",
	1939 => "0000000000000000",1940 => "0000000000000000",1941 => "0000000000000000",
	1942 => "0000000000000000",1943 => "0000000000000000",1944 => "0000000000000000",
	1945 => "0000000000000000",1946 => "0000000000000000",1947 => "0000000000000000",
	1948 => "0000000000000000",1949 => "0000000000000000",1950 => "0000000000000000",
	1951 => "0000000000000000",1952 => "0000000000000000",1953 => "0000000000000000",
	1954 => "0000000000000000",1955 => "0000000000000000",1956 => "0000000000000000",
	1957 => "0000000000000000",1958 => "0000000000000000",1959 => "0000000000000000",
	1960 => "0000000000000000",1961 => "0000000000000000",1962 => "0000000000000000",
	1963 => "0000000000000000",1964 => "0000000000000000",1965 => "0000000000000000",
	1966 => "0000000000000000",1967 => "0000000000000000",1968 => "0000000000000000",
	1969 => "0000000000000000",1970 => "0000000000000000",1971 => "0000000000000000",
	1972 => "0000000000000000",1973 => "0000000000000000",1974 => "0000000000000000",
	1975 => "0000000000000000",1976 => "0000000000000000",1977 => "0000000000000000",
	1978 => "0000000000000000",1979 => "0000000000000000",1980 => "0000000000000000",
	1981 => "0000000000000000",1982 => "0000000000000000",1983 => "0000000000000000",
	1984 => "0000000000000000",1985 => "0000000000000000",1986 => "0000000000000000",
	1987 => "0000000000000000",1988 => "0000000000000000",1989 => "0000000000000000",
	1990 => "0000000000000000",1991 => "0000000000000000",1992 => "0000000000000000",
	1993 => "0000000000000000",1994 => "0000000000000000",1995 => "0000000000000000",
	1996 => "0000000000000000",1997 => "0000000000000000",1998 => "0000000000000000",
	1999 => "0000000000000000",2000 => "0000000000000000",2001 => "0000000000000000",
	2002 => "0000000000000000",2003 => "0000000000000000",2004 => "0000000000000000",
	2005 => "0000000000000000",2006 => "0000000000000000",2007 => "0000000000000000",
	2008 => "0000000000000000",2009 => "0000000000000000",2010 => "0000000000000000",
	2011 => "0000000000000000",2012 => "0000000000000000",2013 => "0000000000000000",
	2014 => "0000000000000000",2015 => "0000000000000000",2016 => "0000000000000000",
	2017 => "0000000000000000",2018 => "0000000000000000",2019 => "0000000000000000",
	2020 => "0000000000000000",2021 => "0000000000000000",2022 => "0000000000000000",
	2023 => "0000000000000000",2024 => "0000000000000000",2025 => "0000000000000000",
	2026 => "0000000000000000",2027 => "0000000000000000",2028 => "0000000000000000",
	2029 => "0000000000000000",2030 => "0000000000000000",2031 => "0000000000000000",
	2032 => "0000000000000000",2033 => "0000000000000000",2034 => "0000000000000000",
	2035 => "0000000000000000",2036 => "0000000000000000",2037 => "0000000000000000",
	2038 => "0000000000000000",2039 => "0000000000000000",2040 => "0000000000000000",
	2041 => "0000000000000000",2042 => "0000000000000000",2043 => "0000000000000000",
	2044 => "0000000000000000",2045 => "0000000000000000",2046 => "0000000000000000",
	2047 => "0000000000000000",2048 => "0000000000000000",2049 => "0000000000000000",
	2050 => "0000000000000000",2051 => "0000000000000000",2052 => "0000000000000000",
	2053 => "0000000000000000",2054 => "0000000000000000",2055 => "0000000000000000",
	2056 => "0000000000000000",2057 => "0000000000000000",2058 => "0000000000000000",
	2059 => "0000000000000000",2060 => "0000000000000000",2061 => "0000000000000000",
	2062 => "0000000000000000",2063 => "0000000000000000",2064 => "0000000000000000",
	2065 => "0000000000000000",2066 => "0000000000000000",2067 => "0000000000000000",
	2068 => "0000000000000000",2069 => "0000000000000000",2070 => "0000000000000000",
	2071 => "0000000000000000",2072 => "0000000000000000",2073 => "0000000000000000",
	2074 => "0000000000000000",2075 => "0000000000000000",2076 => "0000000000000000",
	2077 => "0000000000000000",2078 => "0000000000000000",2079 => "0000000000000000",
	2080 => "0000000000000000",2081 => "0000000000000000",2082 => "0000000000000000",
	2083 => "0000000000000000",2084 => "0000000000000000",2085 => "0000000000000000",
	2086 => "0000000000000000",2087 => "0000000000000000",2088 => "0000000000000000",
	2089 => "0000000000000000",2090 => "0000000000000000",2091 => "0000000000000000",
	2092 => "0000000000000000",2093 => "0000000000000000",2094 => "0000000000000000",
	2095 => "0000000000000000",2096 => "0000000000000000",2097 => "0000000000000000",
	2098 => "0000000000000000",2099 => "0000000000000000",2100 => "0000000000000000",
	2101 => "0000000000000000",2102 => "0000000000000000",2103 => "0000000000000000",
	2104 => "0000000000000000",2105 => "0000000000000000",2106 => "0000000000000000",
	2107 => "0000000000000000",2108 => "0000000000000000",2109 => "0000000000000000",
	2110 => "0000000000000000",2111 => "0000000000000000",2112 => "0000000000000000",
	2113 => "0000000000000000",2114 => "0000000000000000",2115 => "0000000000000000",
	2116 => "0000000000000000",2117 => "0000000000000000",2118 => "0000000000000000",
	2119 => "0000000000000000",2120 => "0000000000000000",2121 => "0000000000000000",
	2122 => "0000000000000000",2123 => "0000000000000000",2124 => "0000000000000000",
	2125 => "0000000000000000",2126 => "0000000000000000",2127 => "0000000000000000",
	2128 => "0000000000000000",2129 => "0000000000000000",2130 => "0000000000000000",
	2131 => "0000000000000000",2132 => "0000000000000000",2133 => "0000000000000000",
	2134 => "0000000000000000",2135 => "0000000000000000",2136 => "0000000000000000",
	2137 => "0000000000000000",2138 => "0000000000000000",2139 => "0000000000000000",
	2140 => "0000000000000000",2141 => "0000000000000000",2142 => "0000000000000000",
	2143 => "0000000000000000",2144 => "0000000000000000",2145 => "0000000000000000",
	2146 => "0000000000000000",2147 => "0000000000000000",2148 => "0000000000000000",
	2149 => "0000000000000000",2150 => "0000000000000000",2151 => "0000000000000000",
	2152 => "0000000000000000",2153 => "0000000000000000",2154 => "0000000000000000",
	2155 => "0000000000000000",2156 => "0000000000000000",2157 => "0000000000000000",
	2158 => "0000000000000000",2159 => "0000000000000000",2160 => "0000000000000000",
	2161 => "0000000000000000",2162 => "0000000000000000",2163 => "0000000000000000",
	2164 => "0000000000000000",2165 => "0000000000000000",2166 => "0000000000000000",
	2167 => "0000000000000000",2168 => "0000000000000000",2169 => "0000000000000000",
	2170 => "0000000000000000",2171 => "0000000000000000",2172 => "0000000000000000",
	2173 => "0000000000000000",2174 => "0000000000000000",2175 => "0000000000000000",
	2176 => "0000000000000000",2177 => "0000000000000000",2178 => "0000000000000000",
	2179 => "0000000000000000",2180 => "0000000000000000",2181 => "0000000000000000",
	2182 => "0000000000000000",2183 => "0000000000000000",2184 => "0000000000000000",
	2185 => "0000000000000000",2186 => "0000000000000000",2187 => "0000000000000000",
	2188 => "0000000000000000",2189 => "0000000000000000",2190 => "0000000000000000",
	2191 => "0000000000000000",2192 => "0000000000000000",2193 => "0000000000000000",
	2194 => "0000000000000000",2195 => "0000000000000000",2196 => "0000000000000000",
	2197 => "0000000000000000",2198 => "0000000000000000",2199 => "0000000000000000",
	2200 => "0000000000000000",2201 => "0000000000000000",2202 => "0000000000000000",
	2203 => "0000000000000000",2204 => "0000000000000000",2205 => "0000000000000000",
	2206 => "0000000000000000",2207 => "0000000000000000",2208 => "0000000000000000",
	2209 => "0000000000000000",2210 => "0000000000000000",2211 => "0000000000000000",
	2212 => "0000000000000000",2213 => "0000000000000000",2214 => "0000000000000000",
	2215 => "0000000000000000",2216 => "0000000000000000",2217 => "0000000000000000",
	2218 => "0000000000000000",2219 => "0000000000000000",2220 => "0000000000000000",
	2221 => "0000000000000000",2222 => "0000000000000000",2223 => "0000000000000000",
	2224 => "0000000000000000",2225 => "0000000000000000",2226 => "0000000000000000",
	2227 => "0000000000000000",2228 => "0000000000000000",2229 => "0000000000000000",
	2230 => "0000000000000000",2231 => "0000000000000000",2232 => "0000000000000000",
	2233 => "0000000000000000",2234 => "0000000000000000",2235 => "0000000000000000",
	2236 => "0000000000000000",2237 => "0000000000000000",2238 => "0000000000000000",
	2239 => "0000000000000000",2240 => "0000000000000000",2241 => "0000000000000000",
	2242 => "0000000000000000",2243 => "0000000000000000",2244 => "0000000000000000",
	2245 => "0000000000000000",2246 => "0000000000000000",2247 => "0000000000000000",
	2248 => "0000000000000000",2249 => "0000000000000000",2250 => "0000000000000000",
	2251 => "0000000000000000",2252 => "0000000000000000",2253 => "0000000000000000",
	2254 => "0000000000000000",2255 => "0000000000000000",2256 => "0000000000000000",
	2257 => "0000000000000000",2258 => "0000000000000000",2259 => "0000000000000000",
	2260 => "0000000000000000",2261 => "0000000000000000",2262 => "0000000000000000",
	2263 => "0000000000000000",2264 => "0000000000000000",2265 => "0000000000000000",
	2266 => "0000000000000000",2267 => "0000000000000000",2268 => "0000000000000000",
	2269 => "0000000000000000",2270 => "0000000000000000",2271 => "0000000000000000",
	2272 => "0000000000000000",2273 => "0000000000000000",2274 => "0000000000000000",
	2275 => "0000000000000000",2276 => "0000000000000000",2277 => "0000000000000000",
	2278 => "0000000000000000",2279 => "0000000000000000",2280 => "0000000000000000",
	2281 => "0000000000000000",2282 => "0000000000000000",2283 => "0000000000000000",
	2284 => "0000000000000000",2285 => "0000000000000000",2286 => "0000000000000000",
	2287 => "0000000000000000",2288 => "0000000000000000",2289 => "0000000000000000",
	2290 => "0000000000000000",2291 => "0000000000000000",2292 => "0000000000000000",
	2293 => "0000000000000000",2294 => "0000000000000000",2295 => "0000000000000000",
	2296 => "0000000000000000",2297 => "0000000000000000",2298 => "0000000000000000",
	2299 => "0000000000000000",2300 => "0000000000000000",2301 => "0000000000000000",
	2302 => "0000000000000000",2303 => "0000000000000000",2304 => "0000000000000000",
	2305 => "0000000000000000",2306 => "0000000000000000",2307 => "0000000000000000",
	2308 => "0000000000000000",2309 => "0000000000000000",2310 => "0000000000000000",
	2311 => "0000000000000000",2312 => "0000000000000000",2313 => "0000000000000000",
	2314 => "0000000000000000",2315 => "0000000000000000",2316 => "0000000000000000",
	2317 => "0000000000000000",2318 => "0000000000000000",2319 => "0000000000000000",
	2320 => "0000000000000000",2321 => "0000000000000000",2322 => "0000000000000000",
	2323 => "0000000000000000",2324 => "0000000000000000",2325 => "0000000000000000",
	2326 => "0000000000000000",2327 => "0000000000000000",2328 => "0000000000000000",
	2329 => "0000000000000000",2330 => "0000000000000000",2331 => "0000000000000000",
	2332 => "0000000000000000",2333 => "0000000000000000",2334 => "0000000000000000",
	2335 => "0000000000000000",2336 => "0000000000000000",2337 => "0000000000000000",
	2338 => "0000000000000000",2339 => "0000000000000000",2340 => "0000000000000000",
	2341 => "0000000000000000",2342 => "0000000000000000",2343 => "0000000000000000",
	2344 => "0000000000000000",2345 => "0000000000000000",2346 => "0000000000000000",
	2347 => "0000000000000000",2348 => "0000000000000000",2349 => "0000000000000000",
	2350 => "0000000000000000",2351 => "0000000000000000",2352 => "0000000000000000",
	2353 => "0000000000000000",2354 => "0000000000000000",2355 => "0000000000000000",
	2356 => "0000000000000000",2357 => "0000000000000000",2358 => "0000000000000000",
	2359 => "0000000000000000",2360 => "0000000000000000",2361 => "0000000000000000",
	2362 => "0000000000000000",2363 => "0000000000000000",2364 => "0000000000000000",
	2365 => "0000000000000000",2366 => "0000000000000000",2367 => "0000000000000000",
	2368 => "0000000000000000",2369 => "0000000000000000",2370 => "0000000000000000",
	2371 => "0000000000000000",2372 => "0000000000000000",2373 => "0000000000000000",
	2374 => "0000000000000000",2375 => "0000000000000000",2376 => "0000000000000000",
	2377 => "0000000000000000",2378 => "0000000000000000",2379 => "0000000000000000",
	2380 => "0000000000000000",2381 => "0000000000000000",2382 => "0000000000000000",
	2383 => "0000000000000000",2384 => "0000000000000000",2385 => "0000000000000000",
	2386 => "0000000000000000",2387 => "0000000000000000",2388 => "0000000000000000",
	2389 => "0000000000000000",2390 => "0000000000000000",2391 => "0000000000000000",
	2392 => "0000000000000000",2393 => "0000000000000000",2394 => "0000000000000000",
	2395 => "0000000000000000",2396 => "0000000000000000",2397 => "0000000000000000",
	2398 => "0000000000000000",2399 => "0000000000000000",2400 => "0000000000000000",
	2401 => "0000000000000000",2402 => "0000000000000000",2403 => "0000000000000000",
	2404 => "0000000000000000",2405 => "0000000000000000",2406 => "0000000000000000",
	2407 => "0000000000000000",2408 => "0000000000000000",2409 => "0000000000000000",
	2410 => "0000000000000000",2411 => "0000000000000000",2412 => "0000000000000000",
	2413 => "0000000000000000",2414 => "0000000000000000",2415 => "0000000000000000",
	2416 => "0000000000000000",2417 => "0000000000000000",2418 => "0000000000000000",
	2419 => "0000000000000000",2420 => "0000000000000000",2421 => "0000000000000000",
	2422 => "0000000000000000",2423 => "0000000000000000",2424 => "0000000000000000",
	2425 => "0000000000000000",2426 => "0000000000000000",2427 => "0000000000000000",
	2428 => "0000000000000000",2429 => "0000000000000000",2430 => "0000000000000000",
	2431 => "0000000000000000",2432 => "0000000000000000",2433 => "0000000000000000",
	2434 => "0000000000000000",2435 => "0000000000000000",2436 => "0000000000000000",
	2437 => "0000000000000000",2438 => "0000000000000000",2439 => "0000000000000000",
	2440 => "0000000000000000",2441 => "0000000000000000",2442 => "0000000000000000",
	2443 => "0000000000000000",2444 => "0000000000000000",2445 => "0000000000000000",
	2446 => "0000000000000000",2447 => "0000000000000000",2448 => "0000000000000000",
	2449 => "0000000000000000",2450 => "0000000000000000",2451 => "0000000000000000",
	2452 => "0000000000000000",2453 => "0000000000000000",2454 => "0000000000000000",
	2455 => "0000000000000000",2456 => "0000000000000000",2457 => "0000000000000000",
	2458 => "0000000000000000",2459 => "0000000000000000",2460 => "0000000000000000",
	2461 => "0000000000000000",2462 => "0000000000000000",2463 => "0000000000000000",
	2464 => "0000000000000000",2465 => "0000000000000000",2466 => "0000000000000000",
	2467 => "0000000000000000",2468 => "0000000000000000",2469 => "0000000000000000",
	2470 => "0000000000000000",2471 => "0000000000000000",2472 => "0000000000000000",
	2473 => "0000000000000000",2474 => "0000000000000000",2475 => "0000000000000000",
	2476 => "0000000000000000",2477 => "0000000000000000",2478 => "0000000000000000",
	2479 => "0000000000000000",2480 => "0000000000000000",2481 => "0000000000000000",
	2482 => "0000000000000000",2483 => "0000000000000000",2484 => "0000000000000000",
	2485 => "0000000000000000",2486 => "0000000000000000",2487 => "0000000000000000",
	2488 => "0000000000000000",2489 => "0000000000000000",2490 => "0000000000000000",
	2491 => "0000000000000000",2492 => "0000000000000000",2493 => "0000000000000000",
	2494 => "0000000000000000",2495 => "0000000000000000",2496 => "0000000000000000",
	2497 => "0000000000000000",2498 => "0000000000000000",2499 => "0000000000000000",
	2500 => "0000000000000000",2501 => "0000000000000000",2502 => "0000000000000000",
	2503 => "0000000000000000",2504 => "0000000000000000",2505 => "0000000000000000",
	2506 => "0000000000000000",2507 => "0000000000000000",2508 => "0000000000000000",
	2509 => "0000000000000000",2510 => "0000000000000000",2511 => "0000000000000000",
	2512 => "0000000000000000",2513 => "0000000000000000",2514 => "0000000000000000",
	2515 => "0000000000000000",2516 => "0000000000000000",2517 => "0000000000000000",
	2518 => "0000000000000000",2519 => "0000000000000000",2520 => "0000000000000000",
	2521 => "0000000000000000",2522 => "0000000000000000",2523 => "0000000000000000",
	2524 => "0000000000000000",2525 => "0000000000000000",2526 => "0000000000000000",
	2527 => "0000000000000000",2528 => "0000000000000000",2529 => "0000000000000000",
	2530 => "0000000000000000",2531 => "0000000000000000",2532 => "0000000000000000",
	2533 => "0000000000000000",2534 => "0000000000000000",2535 => "0000000000000000",
	2536 => "0000000000000000",2537 => "0000000000000000",2538 => "0000000000000000",
	2539 => "0000000000000000",2540 => "0000000000000000",2541 => "0000000000000000",
	2542 => "0000000000000000",2543 => "0000000000000000",2544 => "0000000000000000",
	2545 => "0000000000000000",2546 => "0000000000000000",2547 => "0000000000000000",
	2548 => "0000000000000000",2549 => "0000000000000000",2550 => "0000000000000000",
	2551 => "0000000000000000",2552 => "0000000000000000",2553 => "0000000000000000",
	2554 => "0000000000000000",2555 => "0000000000000000",2556 => "0000000000000000",
	2557 => "0000000000000000",2558 => "0000000000000000",2559 => "0000000000000000",
	2560 => "0000000000000000",2561 => "0000000000000000",2562 => "0000000000000000",
	2563 => "0000000000000000",2564 => "0000000000000000",2565 => "0000000000000000",
	2566 => "0000000000000000",2567 => "0000000000000000",2568 => "0000000000000000",
	2569 => "0000000000000000",2570 => "0000000000000000",2571 => "0000000000000000",
	2572 => "0000000000000000",2573 => "0000000000000000",2574 => "0000000000000000",
	2575 => "0000000000000000",2576 => "0000000000000000",2577 => "0000000000000000",
	2578 => "0000000000000000",2579 => "0000000000000000",2580 => "0000000000000000",
	2581 => "0000000000000000",2582 => "0000000000000000",2583 => "0000000000000000",
	2584 => "0000000000000000",2585 => "0000000000000000",2586 => "0000000000000000",
	2587 => "0000000000000000",2588 => "0000000000000000",2589 => "0000000000000000",
	2590 => "0000000000000000",2591 => "0000000000000000",2592 => "0000000000000000",
	2593 => "0000000000000000",2594 => "0000000000000000",2595 => "0000000000000000",
	2596 => "0000000000000000",2597 => "0000000000000000",2598 => "0000000000000000",
	2599 => "0000000000000000",2600 => "0000000000000000",2601 => "0000000000000000",
	2602 => "0000000000000000",2603 => "0000000000000000",2604 => "0000000000000000",
	2605 => "0000000000000000",2606 => "0000000000000000",2607 => "0000000000000000",
	2608 => "0000000000000000",2609 => "0000000000000000",2610 => "0000000000000000",
	2611 => "0000000000000000",2612 => "0000000000000000",2613 => "0000000000000000",
	2614 => "0000000000000000",2615 => "0000000000000000",2616 => "0000000000000000",
	2617 => "0000000000000000",2618 => "0000000000000000",2619 => "0000000000000000",
	2620 => "0000000000000000",2621 => "0000000000000000",2622 => "0000000000000000",
	2623 => "0000000000000000",2624 => "0000000000000000",2625 => "0000000000000000",
	2626 => "0000000000000000",2627 => "0000000000000000",2628 => "0000000000000000",
	2629 => "0000000000000000",2630 => "0000000000000000",2631 => "0000000000000000",
	2632 => "0000000000000000",2633 => "0000000000000000",2634 => "0000000000000000",
	2635 => "0000000000000000",2636 => "0000000000000000",2637 => "0000000000000000",
	2638 => "0000000000000000",2639 => "0000000000000000",2640 => "0000000000000000",
	2641 => "0000000000000000",2642 => "0000000000000000",2643 => "0000000000000000",
	2644 => "0000000000000000",2645 => "0000000000000000",2646 => "0000000000000000",
	2647 => "0000000000000000",2648 => "0000000000000000",2649 => "0000000000000000",
	2650 => "0000000000000000",2651 => "0000000000000000",2652 => "0000000000000000",
	2653 => "0000000000000000",2654 => "0000000000000000",2655 => "0000000000000000",
	2656 => "0000000000000000",2657 => "0000000000000000",2658 => "0000000000000000",
	2659 => "0000000000000000",2660 => "0000000000000000",2661 => "0000000000000000",
	2662 => "0000000000000000",2663 => "0000000000000000",2664 => "0000000000000000",
	2665 => "0000000000000000",2666 => "0000000000000000",2667 => "0000000000000000",
	2668 => "0000000000000000",2669 => "0000000000000000",2670 => "0000000000000000",
	2671 => "0000000000000000",2672 => "0000000000000000",2673 => "0000000000000000",
	2674 => "0000000000000000",2675 => "0000000000000000",2676 => "0000000000000000",
	2677 => "0000000000000000",2678 => "0000000000000000",2679 => "0000000000000000",
	2680 => "0000000000000000",2681 => "0000000000000000",2682 => "0000000000000000",
	2683 => "0000000000000000",2684 => "0000000000000000",2685 => "0000000000000000",
	2686 => "0000000000000000",2687 => "0000000000000000",2688 => "0000000000000000",
	2689 => "0000000000000000",2690 => "0000000000000000",2691 => "0000000000000000",
	2692 => "0000000000000000",2693 => "0000000000000000",2694 => "0000000000000000",
	2695 => "0000000000000000",2696 => "0000000000000000",2697 => "0000000000000000",
	2698 => "0000000000000000",2699 => "0000000000000000",2700 => "0000000000000000",
	2701 => "0000000000000000",2702 => "0000000000000000",2703 => "0000000000000000",
	2704 => "0000000000000000",2705 => "0000000000000000",2706 => "0000000000000000",
	2707 => "0000000000000000",2708 => "0000000000000000",2709 => "0000000000000000",
	2710 => "0000000000000000",2711 => "0000000000000000",2712 => "0000000000000000",
	2713 => "0000000000000000",2714 => "0000000000000000",2715 => "0000000000000000",
	2716 => "0000000000000000",2717 => "0000000000000000",2718 => "0000000000000000",
	2719 => "0000000000000000",2720 => "0000000000000000",2721 => "0000000000000000",
	2722 => "0000000000000000",2723 => "0000000000000000",2724 => "0000000000000000",
	2725 => "0000000000000000",2726 => "0000000000000000",2727 => "0000000000000000",
	2728 => "0000000000000000",2729 => "0000000000000000",2730 => "0000000000000000",
	2731 => "0000000000000000",2732 => "0000000000000000",2733 => "0000000000000000",
	2734 => "0000000000000000",2735 => "0000000000000000",2736 => "0000000000000000",
	2737 => "0000000000000000",2738 => "0000000000000000",2739 => "0000000000000000",
	2740 => "0000000000000000",2741 => "0000000000000000",2742 => "0000000000000000",
	2743 => "0000000000000000",2744 => "0000000000000000",2745 => "0000000000000000",
	2746 => "0000000000000000",2747 => "0000000000000000",2748 => "0000000000000000",
	2749 => "0000000000000000",2750 => "0000000000000000",2751 => "0000000000000000",
	2752 => "0000000000000000",2753 => "0000000000000000",2754 => "0000000000000000",
	2755 => "0000000000000000",2756 => "0000000000000000",2757 => "0000000000000000",
	2758 => "0000000000000000",2759 => "0000000000000000",2760 => "0000000000000000",
	2761 => "0000000000000000",2762 => "0000000000000000",2763 => "0000000000000000",
	2764 => "0000000000000000",2765 => "0000000000000000",2766 => "0000000000000000",
	2767 => "0000000000000000",2768 => "0000000000000000",2769 => "0000000000000000",
	2770 => "0000000000000000",2771 => "0000000000000000",2772 => "0000000000000000",
	2773 => "0000000000000000",2774 => "0000000000000000",2775 => "0000000000000000",
	2776 => "0000000000000000",2777 => "0000000000000000",2778 => "0000000000000000",
	2779 => "0000000000000000",2780 => "0000000000000000",2781 => "0000000000000000",
	2782 => "0000000000000000",2783 => "0000000000000000",2784 => "0000000000000000",
	2785 => "0000000000000000",2786 => "0000000000000000",2787 => "0000000000000000",
	2788 => "0000000000000000",2789 => "0000000000000000",2790 => "0000000000000000",
	2791 => "0000000000000000",2792 => "0000000000000000",2793 => "0000000000000000",
	2794 => "0000000000000000",2795 => "0000000000000000",2796 => "0000000000000000",
	2797 => "0000000000000000",2798 => "0000000000000000",2799 => "0000000000000000",
	2800 => "0000000000000000",2801 => "0000000000000000",2802 => "0000000000000000",
	2803 => "0000000000000000",2804 => "0000000000000000",2805 => "0000000000000000",
	2806 => "0000000000000000",2807 => "0000000000000000",2808 => "0000000000000000",
	2809 => "0000000000000000",2810 => "0000000000000000",2811 => "0000000000000000",
	2812 => "0000000000000000",2813 => "0000000000000000",2814 => "0000000000000000",
	2815 => "0000000000000000",2816 => "0000000000000000",2817 => "0000000000000000",
	2818 => "0000000000000000",2819 => "0000000000000000",2820 => "0000000000000000",
	2821 => "0000000000000000",2822 => "0000000000000000",2823 => "0000000000000000",
	2824 => "0000000000000000",2825 => "0000000000000000",2826 => "0000000000000000",
	2827 => "0000000000000000",2828 => "0000000000000000",2829 => "0000000000000000",
	2830 => "0000000000000000",2831 => "0000000000000000",2832 => "0000000000000000",
	2833 => "0000000000000000",2834 => "0000000000000000",2835 => "0000000000000000",
	2836 => "0000000000000000",2837 => "0000000000000000",2838 => "0000000000000000",
	2839 => "0000000000000000",2840 => "0000000000000000",2841 => "0000000000000000",
	2842 => "0000000000000000",2843 => "0000000000000000",2844 => "0000000000000000",
	2845 => "0000000000000000",2846 => "0000000000000000",2847 => "0000000000000000",
	2848 => "0000000000000000",2849 => "0000000000000000",2850 => "0000000000000000",
	2851 => "0000000000000000",2852 => "0000000000000000",2853 => "0000000000000000",
	2854 => "0000000000000000",2855 => "0000000000000000",2856 => "0000000000000000",
	2857 => "0000000000000000",2858 => "0000000000000000",2859 => "0000000000000000",
	2860 => "0000000000000000",2861 => "0000000000000000",2862 => "0000000000000000",
	2863 => "0000000000000000",2864 => "0000000000000000",2865 => "0000000000000000",
	2866 => "0000000000000000",2867 => "0000000000000000",2868 => "0000000000000000",
	2869 => "0000000000000000",2870 => "0000000000000000",2871 => "0000000000000000",
	2872 => "0000000000000000",2873 => "0000000000000000",2874 => "0000000000000000",
	2875 => "0000000000000000",2876 => "0000000000000000",2877 => "0000000000000000",
	2878 => "0000000000000000",2879 => "0000000000000000",2880 => "0000000000000000",
	2881 => "0000000000000000",2882 => "0000000000000000",2883 => "0000000000000000",
	2884 => "0000000000000000",2885 => "0000000000000000",2886 => "0000000000000000",
	2887 => "0000000000000000",2888 => "0000000000000000",2889 => "0000000000000000",
	2890 => "0000000000000000",2891 => "0000000000000000",2892 => "0000000000000000",
	2893 => "0000000000000000",2894 => "0000000000000000",2895 => "0000000000000000",
	2896 => "0000000000000000",2897 => "0000000000000000",2898 => "0000000000000000",
	2899 => "0000000000000000",2900 => "0000000000000000",2901 => "0000000000000000",
	2902 => "0000000000000000",2903 => "0000000000000000",2904 => "0000000000000000",
	2905 => "0000000000000000",2906 => "0000000000000000",2907 => "0000000000000000",
	2908 => "0000000000000000",2909 => "0000000000000000",2910 => "0000000000000000",
	2911 => "0000000000000000",2912 => "0000000000000000",2913 => "0000000000000000",
	2914 => "0000000000000000",2915 => "0000000000000000",2916 => "0000000000000000",
	2917 => "0000000000000000",2918 => "0000000000000000",2919 => "0000000000000000",
	2920 => "0000000000000000",2921 => "0000000000000000",2922 => "0000000000000000",
	2923 => "0000000000000000",2924 => "0000000000000000",2925 => "0000000000000000",
	2926 => "0000000000000000",2927 => "0000000000000000",2928 => "0000000000000000",
	2929 => "0000000000000000",2930 => "0000000000000000",2931 => "0000000000000000",
	2932 => "0000000000000000",2933 => "0000000000000000",2934 => "0000000000000000",
	2935 => "0000000000000000",2936 => "0000000000000000",2937 => "0000000000000000",
	2938 => "0000000000000000",2939 => "0000000000000000",2940 => "0000000000000000",
	2941 => "0000000000000000",2942 => "0000000000000000",2943 => "0000000000000000",
	2944 => "0000000000000000",2945 => "0000000000000000",2946 => "0000000000000000",
	2947 => "0000000000000000",2948 => "0000000000000000",2949 => "0000000000000000",
	2950 => "0000000000000000",2951 => "0000000000000000",2952 => "0000000000000000",
	2953 => "0000000000000000",2954 => "0000000000000000",2955 => "0000000000000000",
	2956 => "0000000000000000",2957 => "0000000000000000",2958 => "0000000000000000",
	2959 => "0000000000000000",2960 => "0000000000000000",2961 => "0000000000000000",
	2962 => "0000000000000000",2963 => "0000000000000000",2964 => "0000000000000000",
	2965 => "0000000000000000",2966 => "0000000000000000",2967 => "0000000000000000",
	2968 => "0000000000000000",2969 => "0000000000000000",2970 => "0000000000000000",
	2971 => "0000000000000000",2972 => "0000000000000000",2973 => "0000000000000000",
	2974 => "0000000000000000",2975 => "0000000000000000",2976 => "0000000000000000",
	2977 => "0000000000000000",2978 => "0000000000000000",2979 => "0000000000000000",
	2980 => "0000000000000000",2981 => "0000000000000000",2982 => "0000000000000000",
	2983 => "0000000000000000",2984 => "0000000000000000",2985 => "0000000000000000",
	2986 => "0000000000000000",2987 => "0000000000000000",2988 => "0000000000000000",
	2989 => "0000000000000000",2990 => "0000000000000000",2991 => "0000000000000000",
	2992 => "0000000000000000",2993 => "0000000000000000",2994 => "0000000000000000",
	2995 => "0000000000000000",2996 => "0000000000000000",2997 => "0000000000000000",
	2998 => "0000000000000000",2999 => "0000000000000000",3000 => "0000000000000000",
	3001 => "0000000000000000",3002 => "0000000000000000",3003 => "0000000000000000",
	3004 => "0000000000000000",3005 => "0000000000000000",3006 => "0000000000000000",
	3007 => "0000000000000000",3008 => "0000000000000000",3009 => "0000000000000000",
	others =>"0000000000000000"
);
constant exp_lut_neg : rom_n := (32768 => "0000000100000000",32769 => "0000000011111111",
	32770 => "0000000011111110",32771 => "0000000011111101",32772 => "0000000011111100",
	32773 => "0000000011111011",32774 => "0000000011111010",32775 => "0000000011111001",
	32776 => "0000000011111000",32777 => "0000000011110111",32778 => "0000000011110110",
	32779 => "0000000011110101",32780 => "0000000011110100",32781 => "0000000011110011",
	32782 => "0000000011110010",32783 => "0000000011110001",32784 => "0000000011110000",
	32785 => "0000000011101111",32786 => "0000000011101110",32787 => "0000000011101101",
	32788 => "0000000011101100",32789 => "0000000011101011",32790 => "0000000011101010",
	32791 => "0000000011101010",32792 => "0000000011101001",32793 => "0000000011101000",
	32794 => "0000000011100111",32795 => "0000000011100110",32796 => "0000000011100101",
	32797 => "0000000011100100",32798 => "0000000011100011",32799 => "0000000011100010",
	32800 => "0000000011100001",32801 => "0000000011100001",32802 => "0000000011100000",
	32803 => "0000000011011111",32804 => "0000000011011110",32805 => "0000000011011101",
	32806 => "0000000011011100",32807 => "0000000011011011",32808 => "0000000011011010",
	32809 => "0000000011011010",32810 => "0000000011011001",32811 => "0000000011011000",
	32812 => "0000000011010111",32813 => "0000000011010110",32814 => "0000000011010101",
	32815 => "0000000011010101",32816 => "0000000011010100",32817 => "0000000011010011",
	32818 => "0000000011010010",32819 => "0000000011010001",32820 => "0000000011010000",
	32821 => "0000000011010000",32822 => "0000000011001111",32823 => "0000000011001110",
	32824 => "0000000011001101",32825 => "0000000011001100",32826 => "0000000011001100",
	32827 => "0000000011001011",32828 => "0000000011001010",32829 => "0000000011001001",
	32830 => "0000000011001000",32831 => "0000000011001000",32832 => "0000000011000111",
	32833 => "0000000011000110",32834 => "0000000011000101",32835 => "0000000011000101",
	32836 => "0000000011000100",32837 => "0000000011000011",32838 => "0000000011000010",
	32839 => "0000000011000001",32840 => "0000000011000001",32841 => "0000000011000000",
	32842 => "0000000010111111",32843 => "0000000010111110",32844 => "0000000010111110",
	32845 => "0000000010111101",32846 => "0000000010111100",32847 => "0000000010111100",
	32848 => "0000000010111011",32849 => "0000000010111010",32850 => "0000000010111001",
	32851 => "0000000010111001",32852 => "0000000010111000",32853 => "0000000010110111",
	32854 => "0000000010110110",32855 => "0000000010110110",32856 => "0000000010110101",
	32857 => "0000000010110100",32858 => "0000000010110100",32859 => "0000000010110011",
	32860 => "0000000010110010",32861 => "0000000010110010",32862 => "0000000010110001",
	32863 => "0000000010110000",32864 => "0000000010101111",32865 => "0000000010101111",
	32866 => "0000000010101110",32867 => "0000000010101101",32868 => "0000000010101101",
	32869 => "0000000010101100",32870 => "0000000010101011",32871 => "0000000010101011",
	32872 => "0000000010101010",32873 => "0000000010101001",32874 => "0000000010101001",
	32875 => "0000000010101000",32876 => "0000000010100111",32877 => "0000000010100111",
	32878 => "0000000010100110",32879 => "0000000010100101",32880 => "0000000010100101",
	32881 => "0000000010100100",32882 => "0000000010100011",32883 => "0000000010100011",
	32884 => "0000000010100010",32885 => "0000000010100010",32886 => "0000000010100001",
	32887 => "0000000010100000",32888 => "0000000010100000",32889 => "0000000010011111",
	32890 => "0000000010011110",32891 => "0000000010011110",32892 => "0000000010011101",
	32893 => "0000000010011101",32894 => "0000000010011100",32895 => "0000000010011011",
	32896 => "0000000010011011",32897 => "0000000010011010",32898 => "0000000010011010",
	32899 => "0000000010011001",32900 => "0000000010011000",32901 => "0000000010011000",
	32902 => "0000000010010111",32903 => "0000000010010111",32904 => "0000000010010110",
	32905 => "0000000010010101",32906 => "0000000010010101",32907 => "0000000010010100",
	32908 => "0000000010010100",32909 => "0000000010010011",32910 => "0000000010010011",
	32911 => "0000000010010010",32912 => "0000000010010001",32913 => "0000000010010001",
	32914 => "0000000010010000",32915 => "0000000010010000",32916 => "0000000010001111",
	32917 => "0000000010001111",32918 => "0000000010001110",32919 => "0000000010001101",
	32920 => "0000000010001101",32921 => "0000000010001100",32922 => "0000000010001100",
	32923 => "0000000010001011",32924 => "0000000010001011",32925 => "0000000010001010",
	32926 => "0000000010001010",32927 => "0000000010001001",32928 => "0000000010001001",
	32929 => "0000000010001000",32930 => "0000000010000111",32931 => "0000000010000111",
	32932 => "0000000010000110",32933 => "0000000010000110",32934 => "0000000010000101",
	32935 => "0000000010000101",32936 => "0000000010000100",32937 => "0000000010000100",
	32938 => "0000000010000011",32939 => "0000000010000011",32940 => "0000000010000010",
	32941 => "0000000010000010",32942 => "0000000010000001",32943 => "0000000010000001",
	32944 => "0000000010000000",32945 => "0000000010000000",32946 => "0000000001111111",
	32947 => "0000000001111111",32948 => "0000000001111110",32949 => "0000000001111110",
	32950 => "0000000001111101",32951 => "0000000001111101",32952 => "0000000001111100",
	32953 => "0000000001111100",32954 => "0000000001111011",32955 => "0000000001111011",
	32956 => "0000000001111010",32957 => "0000000001111010",32958 => "0000000001111001",
	32959 => "0000000001111001",32960 => "0000000001111000",32961 => "0000000001111000",
	32962 => "0000000001110111",32963 => "0000000001110111",32964 => "0000000001110111",
	32965 => "0000000001110110",32966 => "0000000001110110",32967 => "0000000001110101",
	32968 => "0000000001110101",32969 => "0000000001110100",32970 => "0000000001110100",
	32971 => "0000000001110011",32972 => "0000000001110011",32973 => "0000000001110010",
	32974 => "0000000001110010",32975 => "0000000001110010",32976 => "0000000001110001",
	32977 => "0000000001110001",32978 => "0000000001110000",32979 => "0000000001110000",
	32980 => "0000000001101111",32981 => "0000000001101111",32982 => "0000000001101110",
	32983 => "0000000001101110",32984 => "0000000001101110",32985 => "0000000001101101",
	32986 => "0000000001101101",32987 => "0000000001101100",32988 => "0000000001101100",
	32989 => "0000000001101011",32990 => "0000000001101011",32991 => "0000000001101011",
	32992 => "0000000001101010",32993 => "0000000001101010",32994 => "0000000001101001",
	32995 => "0000000001101001",32996 => "0000000001101001",32997 => "0000000001101000",
	32998 => "0000000001101000",32999 => "0000000001100111",33000 => "0000000001100111",
	33001 => "0000000001100111",33002 => "0000000001100110",33003 => "0000000001100110",
	33004 => "0000000001100101",33005 => "0000000001100101",33006 => "0000000001100101",
	33007 => "0000000001100100",33008 => "0000000001100100",33009 => "0000000001100011",
	33010 => "0000000001100011",33011 => "0000000001100011",33012 => "0000000001100010",
	33013 => "0000000001100010",33014 => "0000000001100001",33015 => "0000000001100001",
	33016 => "0000000001100001",33017 => "0000000001100000",33018 => "0000000001100000",
	33019 => "0000000001100000",33020 => "0000000001011111",33021 => "0000000001011111",
	33022 => "0000000001011110",33023 => "0000000001011110",33024 => "0000000001011110",
	33025 => "0000000001011101",33026 => "0000000001011101",33027 => "0000000001011101",
	33028 => "0000000001011100",33029 => "0000000001011100",33030 => "0000000001011011",
	33031 => "0000000001011011",33032 => "0000000001011011",33033 => "0000000001011010",
	33034 => "0000000001011010",33035 => "0000000001011010",33036 => "0000000001011001",
	33037 => "0000000001011001",33038 => "0000000001011001",33039 => "0000000001011000",
	33040 => "0000000001011000",33041 => "0000000001011000",33042 => "0000000001010111",
	33043 => "0000000001010111",33044 => "0000000001010111",33045 => "0000000001010110",
	33046 => "0000000001010110",33047 => "0000000001010110",33048 => "0000000001010101",
	33049 => "0000000001010101",33050 => "0000000001010101",33051 => "0000000001010100",
	33052 => "0000000001010100",33053 => "0000000001010100",33054 => "0000000001010011",
	33055 => "0000000001010011",33056 => "0000000001010011",33057 => "0000000001010010",
	33058 => "0000000001010010",33059 => "0000000001010010",33060 => "0000000001010001",
	33061 => "0000000001010001",33062 => "0000000001010001",33063 => "0000000001010000",
	33064 => "0000000001010000",33065 => "0000000001010000",33066 => "0000000001001111",
	33067 => "0000000001001111",33068 => "0000000001001111",33069 => "0000000001001110",
	33070 => "0000000001001110",33071 => "0000000001001110",33072 => "0000000001001110",
	33073 => "0000000001001101",33074 => "0000000001001101",33075 => "0000000001001101",
	33076 => "0000000001001100",33077 => "0000000001001100",33078 => "0000000001001100",
	33079 => "0000000001001011",33080 => "0000000001001011",33081 => "0000000001001011",
	33082 => "0000000001001011",33083 => "0000000001001010",33084 => "0000000001001010",
	33085 => "0000000001001010",33086 => "0000000001001001",33087 => "0000000001001001",
	33088 => "0000000001001001",33089 => "0000000001001001",33090 => "0000000001001000",
	33091 => "0000000001001000",33092 => "0000000001001000",33093 => "0000000001000111",
	33094 => "0000000001000111",33095 => "0000000001000111",33096 => "0000000001000111",
	33097 => "0000000001000110",33098 => "0000000001000110",33099 => "0000000001000110",
	33100 => "0000000001000101",33101 => "0000000001000101",33102 => "0000000001000101",
	33103 => "0000000001000101",33104 => "0000000001000100",33105 => "0000000001000100",
	33106 => "0000000001000100",33107 => "0000000001000100",33108 => "0000000001000011",
	33109 => "0000000001000011",33110 => "0000000001000011",33111 => "0000000001000011",
	33112 => "0000000001000010",33113 => "0000000001000010",33114 => "0000000001000010",
	33115 => "0000000001000010",33116 => "0000000001000001",33117 => "0000000001000001",
	33118 => "0000000001000001",33119 => "0000000001000000",33120 => "0000000001000000",
	33121 => "0000000001000000",33122 => "0000000001000000",33123 => "0000000000111111",
	33124 => "0000000000111111",33125 => "0000000000111111",33126 => "0000000000111111",
	33127 => "0000000000111110",33128 => "0000000000111110",33129 => "0000000000111110",
	33130 => "0000000000111110",33131 => "0000000000111110",33132 => "0000000000111101",
	33133 => "0000000000111101",33134 => "0000000000111101",33135 => "0000000000111101",
	33136 => "0000000000111100",33137 => "0000000000111100",33138 => "0000000000111100",
	33139 => "0000000000111100",33140 => "0000000000111011",33141 => "0000000000111011",
	33142 => "0000000000111011",33143 => "0000000000111011",33144 => "0000000000111010",
	33145 => "0000000000111010",33146 => "0000000000111010",33147 => "0000000000111010",
	33148 => "0000000000111010",33149 => "0000000000111001",33150 => "0000000000111001",
	33151 => "0000000000111001",33152 => "0000000000111001",33153 => "0000000000111000",
	33154 => "0000000000111000",33155 => "0000000000111000",33156 => "0000000000111000",
	33157 => "0000000000111000",33158 => "0000000000110111",33159 => "0000000000110111",
	33160 => "0000000000110111",33161 => "0000000000110111",33162 => "0000000000110110",
	33163 => "0000000000110110",33164 => "0000000000110110",33165 => "0000000000110110",
	33166 => "0000000000110110",33167 => "0000000000110101",33168 => "0000000000110101",
	33169 => "0000000000110101",33170 => "0000000000110101",33171 => "0000000000110101",
	33172 => "0000000000110100",33173 => "0000000000110100",33174 => "0000000000110100",
	33175 => "0000000000110100",33176 => "0000000000110100",33177 => "0000000000110011",
	33178 => "0000000000110011",33179 => "0000000000110011",33180 => "0000000000110011",
	33181 => "0000000000110011",33182 => "0000000000110010",33183 => "0000000000110010",
	33184 => "0000000000110010",33185 => "0000000000110010",33186 => "0000000000110010",
	33187 => "0000000000110001",33188 => "0000000000110001",33189 => "0000000000110001",
	33190 => "0000000000110001",33191 => "0000000000110001",33192 => "0000000000110000",
	33193 => "0000000000110000",33194 => "0000000000110000",33195 => "0000000000110000",
	33196 => "0000000000110000",33197 => "0000000000101111",33198 => "0000000000101111",
	33199 => "0000000000101111",33200 => "0000000000101111",33201 => "0000000000101111",
	33202 => "0000000000101110",33203 => "0000000000101110",33204 => "0000000000101110",
	33205 => "0000000000101110",33206 => "0000000000101110",33207 => "0000000000101110",
	33208 => "0000000000101101",33209 => "0000000000101101",33210 => "0000000000101101",
	33211 => "0000000000101101",33212 => "0000000000101101",33213 => "0000000000101101",
	33214 => "0000000000101100",33215 => "0000000000101100",33216 => "0000000000101100",
	33217 => "0000000000101100",33218 => "0000000000101100",33219 => "0000000000101011",
	33220 => "0000000000101011",33221 => "0000000000101011",33222 => "0000000000101011",
	33223 => "0000000000101011",33224 => "0000000000101011",33225 => "0000000000101010",
	33226 => "0000000000101010",33227 => "0000000000101010",33228 => "0000000000101010",
	33229 => "0000000000101010",33230 => "0000000000101010",33231 => "0000000000101001",
	33232 => "0000000000101001",33233 => "0000000000101001",33234 => "0000000000101001",
	33235 => "0000000000101001",33236 => "0000000000101001",33237 => "0000000000101000",
	33238 => "0000000000101000",33239 => "0000000000101000",33240 => "0000000000101000",
	33241 => "0000000000101000",33242 => "0000000000101000",33243 => "0000000000101000",
	33244 => "0000000000100111",33245 => "0000000000100111",33246 => "0000000000100111",
	33247 => "0000000000100111",33248 => "0000000000100111",33249 => "0000000000100111",
	33250 => "0000000000100110",33251 => "0000000000100110",33252 => "0000000000100110",
	33253 => "0000000000100110",33254 => "0000000000100110",33255 => "0000000000100110",
	33256 => "0000000000100110",33257 => "0000000000100101",33258 => "0000000000100101",
	33259 => "0000000000100101",33260 => "0000000000100101",33261 => "0000000000100101",
	33262 => "0000000000100101",33263 => "0000000000100101",33264 => "0000000000100100",
	33265 => "0000000000100100",33266 => "0000000000100100",33267 => "0000000000100100",
	33268 => "0000000000100100",33269 => "0000000000100100",33270 => "0000000000100100",
	33271 => "0000000000100011",33272 => "0000000000100011",33273 => "0000000000100011",
	33274 => "0000000000100011",33275 => "0000000000100011",33276 => "0000000000100011",
	33277 => "0000000000100011",33278 => "0000000000100010",33279 => "0000000000100010",
	33280 => "0000000000100010",33281 => "0000000000100010",33282 => "0000000000100010",
	33283 => "0000000000100010",33284 => "0000000000100010",33285 => "0000000000100001",
	33286 => "0000000000100001",33287 => "0000000000100001",33288 => "0000000000100001",
	33289 => "0000000000100001",33290 => "0000000000100001",33291 => "0000000000100001",
	33292 => "0000000000100001",33293 => "0000000000100000",33294 => "0000000000100000",
	33295 => "0000000000100000",33296 => "0000000000100000",33297 => "0000000000100000",
	33298 => "0000000000100000",33299 => "0000000000100000",33300 => "0000000000100000",
	33301 => "0000000000011111",33302 => "0000000000011111",33303 => "0000000000011111",
	33304 => "0000000000011111",33305 => "0000000000011111",33306 => "0000000000011111",
	33307 => "0000000000011111",33308 => "0000000000011111",33309 => "0000000000011110",
	33310 => "0000000000011110",33311 => "0000000000011110",33312 => "0000000000011110",
	33313 => "0000000000011110",33314 => "0000000000011110",33315 => "0000000000011110",
	33316 => "0000000000011110",33317 => "0000000000011101",33318 => "0000000000011101",
	33319 => "0000000000011101",33320 => "0000000000011101",33321 => "0000000000011101",
	33322 => "0000000000011101",33323 => "0000000000011101",33324 => "0000000000011101",
	33325 => "0000000000011101",33326 => "0000000000011100",33327 => "0000000000011100",
	33328 => "0000000000011100",33329 => "0000000000011100",33330 => "0000000000011100",
	33331 => "0000000000011100",33332 => "0000000000011100",33333 => "0000000000011100",
	33334 => "0000000000011100",33335 => "0000000000011011",33336 => "0000000000011011",
	33337 => "0000000000011011",33338 => "0000000000011011",33339 => "0000000000011011",
	33340 => "0000000000011011",33341 => "0000000000011011",33342 => "0000000000011011",
	33343 => "0000000000011011",33344 => "0000000000011010",33345 => "0000000000011010",
	33346 => "0000000000011010",33347 => "0000000000011010",33348 => "0000000000011010",
	33349 => "0000000000011010",33350 => "0000000000011010",33351 => "0000000000011010",
	33352 => "0000000000011010",33353 => "0000000000011010",33354 => "0000000000011001",
	33355 => "0000000000011001",33356 => "0000000000011001",33357 => "0000000000011001",
	33358 => "0000000000011001",33359 => "0000000000011001",33360 => "0000000000011001",
	33361 => "0000000000011001",33362 => "0000000000011001",33363 => "0000000000011001",
	33364 => "0000000000011000",33365 => "0000000000011000",33366 => "0000000000011000",
	33367 => "0000000000011000",33368 => "0000000000011000",33369 => "0000000000011000",
	33370 => "0000000000011000",33371 => "0000000000011000",33372 => "0000000000011000",
	33373 => "0000000000011000",33374 => "0000000000010111",33375 => "0000000000010111",
	33376 => "0000000000010111",33377 => "0000000000010111",33378 => "0000000000010111",
	33379 => "0000000000010111",33380 => "0000000000010111",33381 => "0000000000010111",
	33382 => "0000000000010111",33383 => "0000000000010111",33384 => "0000000000010111",
	33385 => "0000000000010110",33386 => "0000000000010110",33387 => "0000000000010110",
	33388 => "0000000000010110",33389 => "0000000000010110",33390 => "0000000000010110",
	33391 => "0000000000010110",33392 => "0000000000010110",33393 => "0000000000010110",
	33394 => "0000000000010110",33395 => "0000000000010110",33396 => "0000000000010110",
	33397 => "0000000000010101",33398 => "0000000000010101",33399 => "0000000000010101",
	33400 => "0000000000010101",33401 => "0000000000010101",33402 => "0000000000010101",
	33403 => "0000000000010101",33404 => "0000000000010101",33405 => "0000000000010101",
	33406 => "0000000000010101",33407 => "0000000000010101",33408 => "0000000000010101",
	33409 => "0000000000010100",33410 => "0000000000010100",33411 => "0000000000010100",
	33412 => "0000000000010100",33413 => "0000000000010100",33414 => "0000000000010100",
	33415 => "0000000000010100",33416 => "0000000000010100",33417 => "0000000000010100",
	33418 => "0000000000010100",33419 => "0000000000010100",33420 => "0000000000010100",
	33421 => "0000000000010011",33422 => "0000000000010011",33423 => "0000000000010011",
	33424 => "0000000000010011",33425 => "0000000000010011",33426 => "0000000000010011",
	33427 => "0000000000010011",33428 => "0000000000010011",33429 => "0000000000010011",
	33430 => "0000000000010011",33431 => "0000000000010011",33432 => "0000000000010011",
	33433 => "0000000000010011",33434 => "0000000000010010",33435 => "0000000000010010",
	33436 => "0000000000010010",33437 => "0000000000010010",33438 => "0000000000010010",
	33439 => "0000000000010010",33440 => "0000000000010010",33441 => "0000000000010010",
	33442 => "0000000000010010",33443 => "0000000000010010",33444 => "0000000000010010",
	33445 => "0000000000010010",33446 => "0000000000010010",33447 => "0000000000010010",
	33448 => "0000000000010001",33449 => "0000000000010001",33450 => "0000000000010001",
	33451 => "0000000000010001",33452 => "0000000000010001",33453 => "0000000000010001",
	33454 => "0000000000010001",33455 => "0000000000010001",33456 => "0000000000010001",
	33457 => "0000000000010001",33458 => "0000000000010001",33459 => "0000000000010001",
	33460 => "0000000000010001",33461 => "0000000000010001",33462 => "0000000000010001",
	33463 => "0000000000010000",33464 => "0000000000010000",33465 => "0000000000010000",
	33466 => "0000000000010000",33467 => "0000000000010000",33468 => "0000000000010000",
	33469 => "0000000000010000",33470 => "0000000000010000",33471 => "0000000000010000",
	33472 => "0000000000010000",33473 => "0000000000010000",33474 => "0000000000010000",
	33475 => "0000000000010000",33476 => "0000000000010000",33477 => "0000000000010000",
	33478 => "0000000000001111",33479 => "0000000000001111",33480 => "0000000000001111",
	33481 => "0000000000001111",33482 => "0000000000001111",33483 => "0000000000001111",
	33484 => "0000000000001111",33485 => "0000000000001111",33486 => "0000000000001111",
	33487 => "0000000000001111",33488 => "0000000000001111",33489 => "0000000000001111",
	33490 => "0000000000001111",33491 => "0000000000001111",33492 => "0000000000001111",
	33493 => "0000000000001111",33494 => "0000000000001111",33495 => "0000000000001110",
	33496 => "0000000000001110",33497 => "0000000000001110",33498 => "0000000000001110",
	33499 => "0000000000001110",33500 => "0000000000001110",33501 => "0000000000001110",
	33502 => "0000000000001110",33503 => "0000000000001110",33504 => "0000000000001110",
	33505 => "0000000000001110",33506 => "0000000000001110",33507 => "0000000000001110",
	33508 => "0000000000001110",33509 => "0000000000001110",33510 => "0000000000001110",
	33511 => "0000000000001110",33512 => "0000000000001101",33513 => "0000000000001101",
	33514 => "0000000000001101",33515 => "0000000000001101",33516 => "0000000000001101",
	33517 => "0000000000001101",33518 => "0000000000001101",33519 => "0000000000001101",
	33520 => "0000000000001101",33521 => "0000000000001101",33522 => "0000000000001101",
	33523 => "0000000000001101",33524 => "0000000000001101",33525 => "0000000000001101",
	33526 => "0000000000001101",33527 => "0000000000001101",33528 => "0000000000001101",
	33529 => "0000000000001101",33530 => "0000000000001101",33531 => "0000000000001100",
	33532 => "0000000000001100",33533 => "0000000000001100",33534 => "0000000000001100",
	33535 => "0000000000001100",33536 => "0000000000001100",33537 => "0000000000001100",
	33538 => "0000000000001100",33539 => "0000000000001100",33540 => "0000000000001100",
	33541 => "0000000000001100",33542 => "0000000000001100",33543 => "0000000000001100",
	33544 => "0000000000001100",33545 => "0000000000001100",33546 => "0000000000001100",
	33547 => "0000000000001100",33548 => "0000000000001100",33549 => "0000000000001100",
	33550 => "0000000000001100",33551 => "0000000000001100",33552 => "0000000000001011",
	33553 => "0000000000001011",33554 => "0000000000001011",33555 => "0000000000001011",
	33556 => "0000000000001011",33557 => "0000000000001011",33558 => "0000000000001011",
	33559 => "0000000000001011",33560 => "0000000000001011",33561 => "0000000000001011",
	33562 => "0000000000001011",33563 => "0000000000001011",33564 => "0000000000001011",
	33565 => "0000000000001011",33566 => "0000000000001011",33567 => "0000000000001011",
	33568 => "0000000000001011",33569 => "0000000000001011",33570 => "0000000000001011",
	33571 => "0000000000001011",33572 => "0000000000001011",33573 => "0000000000001011",
	33574 => "0000000000001010",33575 => "0000000000001010",33576 => "0000000000001010",
	33577 => "0000000000001010",33578 => "0000000000001010",33579 => "0000000000001010",
	33580 => "0000000000001010",33581 => "0000000000001010",33582 => "0000000000001010",
	33583 => "0000000000001010",33584 => "0000000000001010",33585 => "0000000000001010",
	33586 => "0000000000001010",33587 => "0000000000001010",33588 => "0000000000001010",
	33589 => "0000000000001010",33590 => "0000000000001010",33591 => "0000000000001010",
	33592 => "0000000000001010",33593 => "0000000000001010",33594 => "0000000000001010",
	33595 => "0000000000001010",33596 => "0000000000001010",33597 => "0000000000001010",
	33598 => "0000000000001010",33599 => "0000000000001001",33600 => "0000000000001001",
	33601 => "0000000000001001",33602 => "0000000000001001",33603 => "0000000000001001",
	33604 => "0000000000001001",33605 => "0000000000001001",33606 => "0000000000001001",
	33607 => "0000000000001001",33608 => "0000000000001001",33609 => "0000000000001001",
	33610 => "0000000000001001",33611 => "0000000000001001",33612 => "0000000000001001",
	33613 => "0000000000001001",33614 => "0000000000001001",33615 => "0000000000001001",
	33616 => "0000000000001001",33617 => "0000000000001001",33618 => "0000000000001001",
	33619 => "0000000000001001",33620 => "0000000000001001",33621 => "0000000000001001",
	33622 => "0000000000001001",33623 => "0000000000001001",33624 => "0000000000001001",
	33625 => "0000000000001001",33626 => "0000000000001000",33627 => "0000000000001000",
	33628 => "0000000000001000",33629 => "0000000000001000",33630 => "0000000000001000",
	33631 => "0000000000001000",33632 => "0000000000001000",33633 => "0000000000001000",
	33634 => "0000000000001000",33635 => "0000000000001000",33636 => "0000000000001000",
	33637 => "0000000000001000",33638 => "0000000000001000",33639 => "0000000000001000",
	33640 => "0000000000001000",33641 => "0000000000001000",33642 => "0000000000001000",
	33643 => "0000000000001000",33644 => "0000000000001000",33645 => "0000000000001000",
	33646 => "0000000000001000",33647 => "0000000000001000",33648 => "0000000000001000",
	33649 => "0000000000001000",33650 => "0000000000001000",33651 => "0000000000001000",
	33652 => "0000000000001000",33653 => "0000000000001000",33654 => "0000000000001000",
	33655 => "0000000000001000",33656 => "0000000000000111",33657 => "0000000000000111",
	33658 => "0000000000000111",33659 => "0000000000000111",33660 => "0000000000000111",
	33661 => "0000000000000111",33662 => "0000000000000111",33663 => "0000000000000111",
	33664 => "0000000000000111",33665 => "0000000000000111",33666 => "0000000000000111",
	33667 => "0000000000000111",33668 => "0000000000000111",33669 => "0000000000000111",
	33670 => "0000000000000111",33671 => "0000000000000111",33672 => "0000000000000111",
	33673 => "0000000000000111",33674 => "0000000000000111",33675 => "0000000000000111",
	33676 => "0000000000000111",33677 => "0000000000000111",33678 => "0000000000000111",
	33679 => "0000000000000111",33680 => "0000000000000111",33681 => "0000000000000111",
	33682 => "0000000000000111",33683 => "0000000000000111",33684 => "0000000000000111",
	33685 => "0000000000000111",33686 => "0000000000000111",33687 => "0000000000000111",
	33688 => "0000000000000111",33689 => "0000000000000111",33690 => "0000000000000110",
	33691 => "0000000000000110",33692 => "0000000000000110",33693 => "0000000000000110",
	33694 => "0000000000000110",33695 => "0000000000000110",33696 => "0000000000000110",
	33697 => "0000000000000110",33698 => "0000000000000110",33699 => "0000000000000110",
	33700 => "0000000000000110",33701 => "0000000000000110",33702 => "0000000000000110",
	33703 => "0000000000000110",33704 => "0000000000000110",33705 => "0000000000000110",
	33706 => "0000000000000110",33707 => "0000000000000110",33708 => "0000000000000110",
	33709 => "0000000000000110",33710 => "0000000000000110",33711 => "0000000000000110",
	33712 => "0000000000000110",33713 => "0000000000000110",33714 => "0000000000000110",
	33715 => "0000000000000110",33716 => "0000000000000110",33717 => "0000000000000110",
	33718 => "0000000000000110",33719 => "0000000000000110",33720 => "0000000000000110",
	33721 => "0000000000000110",33722 => "0000000000000110",33723 => "0000000000000110",
	33724 => "0000000000000110",33725 => "0000000000000110",33726 => "0000000000000110",
	33727 => "0000000000000110",33728 => "0000000000000110",33729 => "0000000000000101",
	33730 => "0000000000000101",33731 => "0000000000000101",33732 => "0000000000000101",
	33733 => "0000000000000101",33734 => "0000000000000101",33735 => "0000000000000101",
	33736 => "0000000000000101",33737 => "0000000000000101",33738 => "0000000000000101",
	33739 => "0000000000000101",33740 => "0000000000000101",33741 => "0000000000000101",
	33742 => "0000000000000101",33743 => "0000000000000101",33744 => "0000000000000101",
	33745 => "0000000000000101",33746 => "0000000000000101",33747 => "0000000000000101",
	33748 => "0000000000000101",33749 => "0000000000000101",33750 => "0000000000000101",
	33751 => "0000000000000101",33752 => "0000000000000101",33753 => "0000000000000101",
	33754 => "0000000000000101",33755 => "0000000000000101",33756 => "0000000000000101",
	33757 => "0000000000000101",33758 => "0000000000000101",33759 => "0000000000000101",
	33760 => "0000000000000101",33761 => "0000000000000101",33762 => "0000000000000101",
	33763 => "0000000000000101",33764 => "0000000000000101",33765 => "0000000000000101",
	33766 => "0000000000000101",33767 => "0000000000000101",33768 => "0000000000000101",
	33769 => "0000000000000101",33770 => "0000000000000101",33771 => "0000000000000101",
	33772 => "0000000000000101",33773 => "0000000000000101",33774 => "0000000000000101",
	33775 => "0000000000000101",33776 => "0000000000000100",33777 => "0000000000000100",
	33778 => "0000000000000100",33779 => "0000000000000100",33780 => "0000000000000100",
	33781 => "0000000000000100",33782 => "0000000000000100",33783 => "0000000000000100",
	33784 => "0000000000000100",33785 => "0000000000000100",33786 => "0000000000000100",
	33787 => "0000000000000100",33788 => "0000000000000100",33789 => "0000000000000100",
	33790 => "0000000000000100",33791 => "0000000000000100",33792 => "0000000000000100",
	33793 => "0000000000000100",33794 => "0000000000000100",33795 => "0000000000000100",
	33796 => "0000000000000100",33797 => "0000000000000100",33798 => "0000000000000100",
	33799 => "0000000000000100",33800 => "0000000000000100",33801 => "0000000000000100",
	33802 => "0000000000000100",33803 => "0000000000000100",33804 => "0000000000000100",
	33805 => "0000000000000100",33806 => "0000000000000100",33807 => "0000000000000100",
	33808 => "0000000000000100",33809 => "0000000000000100",33810 => "0000000000000100",
	33811 => "0000000000000100",33812 => "0000000000000100",33813 => "0000000000000100",
	33814 => "0000000000000100",33815 => "0000000000000100",33816 => "0000000000000100",
	33817 => "0000000000000100",33818 => "0000000000000100",33819 => "0000000000000100",
	33820 => "0000000000000100",33821 => "0000000000000100",33822 => "0000000000000100",
	33823 => "0000000000000100",33824 => "0000000000000100",33825 => "0000000000000100",
	33826 => "0000000000000100",33827 => "0000000000000100",33828 => "0000000000000100",
	33829 => "0000000000000100",33830 => "0000000000000100",33831 => "0000000000000100",
	33832 => "0000000000000100",33833 => "0000000000000011",33834 => "0000000000000011",
	33835 => "0000000000000011",33836 => "0000000000000011",33837 => "0000000000000011",
	33838 => "0000000000000011",33839 => "0000000000000011",33840 => "0000000000000011",
	33841 => "0000000000000011",33842 => "0000000000000011",33843 => "0000000000000011",
	33844 => "0000000000000011",33845 => "0000000000000011",33846 => "0000000000000011",
	33847 => "0000000000000011",33848 => "0000000000000011",33849 => "0000000000000011",
	33850 => "0000000000000011",33851 => "0000000000000011",33852 => "0000000000000011",
	33853 => "0000000000000011",33854 => "0000000000000011",33855 => "0000000000000011",
	33856 => "0000000000000011",33857 => "0000000000000011",33858 => "0000000000000011",
	33859 => "0000000000000011",33860 => "0000000000000011",33861 => "0000000000000011",
	33862 => "0000000000000011",33863 => "0000000000000011",33864 => "0000000000000011",
	33865 => "0000000000000011",33866 => "0000000000000011",33867 => "0000000000000011",
	33868 => "0000000000000011",33869 => "0000000000000011",33870 => "0000000000000011",
	33871 => "0000000000000011",33872 => "0000000000000011",33873 => "0000000000000011",
	33874 => "0000000000000011",33875 => "0000000000000011",33876 => "0000000000000011",
	33877 => "0000000000000011",33878 => "0000000000000011",33879 => "0000000000000011",
	33880 => "0000000000000011",33881 => "0000000000000011",33882 => "0000000000000011",
	33883 => "0000000000000011",33884 => "0000000000000011",33885 => "0000000000000011",
	33886 => "0000000000000011",33887 => "0000000000000011",33888 => "0000000000000011",
	33889 => "0000000000000011",33890 => "0000000000000011",33891 => "0000000000000011",
	33892 => "0000000000000011",33893 => "0000000000000011",33894 => "0000000000000011",
	33895 => "0000000000000011",33896 => "0000000000000011",33897 => "0000000000000011",
	33898 => "0000000000000011",33899 => "0000000000000011",33900 => "0000000000000011",
	33901 => "0000000000000011",33902 => "0000000000000011",33903 => "0000000000000011",
	33904 => "0000000000000011",33905 => "0000000000000011",33906 => "0000000000000011",
	33907 => "0000000000000010",33908 => "0000000000000010",33909 => "0000000000000010",
	33910 => "0000000000000010",33911 => "0000000000000010",33912 => "0000000000000010",
	33913 => "0000000000000010",33914 => "0000000000000010",33915 => "0000000000000010",
	33916 => "0000000000000010",33917 => "0000000000000010",33918 => "0000000000000010",
	33919 => "0000000000000010",33920 => "0000000000000010",33921 => "0000000000000010",
	33922 => "0000000000000010",33923 => "0000000000000010",33924 => "0000000000000010",
	33925 => "0000000000000010",33926 => "0000000000000010",33927 => "0000000000000010",
	33928 => "0000000000000010",33929 => "0000000000000010",33930 => "0000000000000010",
	33931 => "0000000000000010",33932 => "0000000000000010",33933 => "0000000000000010",
	33934 => "0000000000000010",33935 => "0000000000000010",33936 => "0000000000000010",
	33937 => "0000000000000010",33938 => "0000000000000010",33939 => "0000000000000010",
	33940 => "0000000000000010",33941 => "0000000000000010",33942 => "0000000000000010",
	33943 => "0000000000000010",33944 => "0000000000000010",33945 => "0000000000000010",
	33946 => "0000000000000010",33947 => "0000000000000010",33948 => "0000000000000010",
	33949 => "0000000000000010",33950 => "0000000000000010",33951 => "0000000000000010",
	33952 => "0000000000000010",33953 => "0000000000000010",33954 => "0000000000000010",
	33955 => "0000000000000010",33956 => "0000000000000010",33957 => "0000000000000010",
	33958 => "0000000000000010",33959 => "0000000000000010",33960 => "0000000000000010",
	33961 => "0000000000000010",33962 => "0000000000000010",33963 => "0000000000000010",
	33964 => "0000000000000010",33965 => "0000000000000010",33966 => "0000000000000010",
	33967 => "0000000000000010",33968 => "0000000000000010",33969 => "0000000000000010",
	33970 => "0000000000000010",33971 => "0000000000000010",33972 => "0000000000000010",
	33973 => "0000000000000010",33974 => "0000000000000010",33975 => "0000000000000010",
	33976 => "0000000000000010",33977 => "0000000000000010",33978 => "0000000000000010",
	33979 => "0000000000000010",33980 => "0000000000000010",33981 => "0000000000000010",
	33982 => "0000000000000010",33983 => "0000000000000010",33984 => "0000000000000010",
	33985 => "0000000000000010",33986 => "0000000000000010",33987 => "0000000000000010",
	33988 => "0000000000000010",33989 => "0000000000000010",33990 => "0000000000000010",
	33991 => "0000000000000010",33992 => "0000000000000010",33993 => "0000000000000010",
	33994 => "0000000000000010",33995 => "0000000000000010",33996 => "0000000000000010",
	33997 => "0000000000000010",33998 => "0000000000000010",33999 => "0000000000000010",
	34000 => "0000000000000010",34001 => "0000000000000010",34002 => "0000000000000010",
	34003 => "0000000000000010",34004 => "0000000000000010",34005 => "0000000000000010",
	34006 => "0000000000000010",34007 => "0000000000000010",34008 => "0000000000000010",
	34009 => "0000000000000010",34010 => "0000000000000010",34011 => "0000000000000001",
	34012 => "0000000000000001",34013 => "0000000000000001",34014 => "0000000000000001",
	34015 => "0000000000000001",34016 => "0000000000000001",34017 => "0000000000000001",
	34018 => "0000000000000001",34019 => "0000000000000001",34020 => "0000000000000001",
	34021 => "0000000000000001",34022 => "0000000000000001",34023 => "0000000000000001",
	34024 => "0000000000000001",34025 => "0000000000000001",34026 => "0000000000000001",
	34027 => "0000000000000001",34028 => "0000000000000001",34029 => "0000000000000001",
	34030 => "0000000000000001",34031 => "0000000000000001",34032 => "0000000000000001",
	34033 => "0000000000000001",34034 => "0000000000000001",34035 => "0000000000000001",
	34036 => "0000000000000001",34037 => "0000000000000001",34038 => "0000000000000001",
	34039 => "0000000000000001",34040 => "0000000000000001",34041 => "0000000000000001",
	34042 => "0000000000000001",34043 => "0000000000000001",34044 => "0000000000000001",
	34045 => "0000000000000001",34046 => "0000000000000001",34047 => "0000000000000001",
	34048 => "0000000000000001",34049 => "0000000000000001",34050 => "0000000000000001",
	34051 => "0000000000000001",34052 => "0000000000000001",34053 => "0000000000000001",
	34054 => "0000000000000001",34055 => "0000000000000001",34056 => "0000000000000001",
	34057 => "0000000000000001",34058 => "0000000000000001",34059 => "0000000000000001",
	34060 => "0000000000000001",34061 => "0000000000000001",34062 => "0000000000000001",
	34063 => "0000000000000001",34064 => "0000000000000001",34065 => "0000000000000001",
	34066 => "0000000000000001",34067 => "0000000000000001",34068 => "0000000000000001",
	34069 => "0000000000000001",34070 => "0000000000000001",34071 => "0000000000000001",
	34072 => "0000000000000001",34073 => "0000000000000001",34074 => "0000000000000001",
	34075 => "0000000000000001",34076 => "0000000000000001",34077 => "0000000000000001",
	34078 => "0000000000000001",34079 => "0000000000000001",34080 => "0000000000000001",
	34081 => "0000000000000001",34082 => "0000000000000001",34083 => "0000000000000001",
	34084 => "0000000000000001",34085 => "0000000000000001",34086 => "0000000000000001",
	34087 => "0000000000000001",34088 => "0000000000000001",34089 => "0000000000000001",
	34090 => "0000000000000001",34091 => "0000000000000001",34092 => "0000000000000001",
	34093 => "0000000000000001",34094 => "0000000000000001",34095 => "0000000000000001",
	34096 => "0000000000000001",34097 => "0000000000000001",34098 => "0000000000000001",
	34099 => "0000000000000001",34100 => "0000000000000001",34101 => "0000000000000001",
	34102 => "0000000000000001",34103 => "0000000000000001",34104 => "0000000000000001",
	34105 => "0000000000000001",34106 => "0000000000000001",34107 => "0000000000000001",
	34108 => "0000000000000001",34109 => "0000000000000001",34110 => "0000000000000001",
	34111 => "0000000000000001",34112 => "0000000000000001",34113 => "0000000000000001",
	34114 => "0000000000000001",34115 => "0000000000000001",34116 => "0000000000000001",
	34117 => "0000000000000001",34118 => "0000000000000001",34119 => "0000000000000001",
	34120 => "0000000000000001",34121 => "0000000000000001",34122 => "0000000000000001",
	34123 => "0000000000000001",34124 => "0000000000000001",34125 => "0000000000000001",
	34126 => "0000000000000001",34127 => "0000000000000001",34128 => "0000000000000001",
	34129 => "0000000000000001",34130 => "0000000000000001",34131 => "0000000000000001",
	34132 => "0000000000000001",34133 => "0000000000000001",34134 => "0000000000000001",
	34135 => "0000000000000001",34136 => "0000000000000001",34137 => "0000000000000001",
	34138 => "0000000000000001",34139 => "0000000000000001",34140 => "0000000000000001",
	34141 => "0000000000000001",34142 => "0000000000000001",34143 => "0000000000000001",
	34144 => "0000000000000001",34145 => "0000000000000001",34146 => "0000000000000001",
	34147 => "0000000000000001",34148 => "0000000000000001",34149 => "0000000000000001",
	34150 => "0000000000000001",34151 => "0000000000000001",34152 => "0000000000000001",
	34153 => "0000000000000001",34154 => "0000000000000001",34155 => "0000000000000001",
	34156 => "0000000000000001",34157 => "0000000000000001",34158 => "0000000000000001",
	34159 => "0000000000000001",34160 => "0000000000000001",34161 => "0000000000000001",
	34162 => "0000000000000001",34163 => "0000000000000001",34164 => "0000000000000001",
	34165 => "0000000000000001",34166 => "0000000000000001",34167 => "0000000000000001",
	34168 => "0000000000000001",34169 => "0000000000000001",34170 => "0000000000000001",
	34171 => "0000000000000001",34172 => "0000000000000001",34173 => "0000000000000001",
	34174 => "0000000000000001",34175 => "0000000000000001",34176 => "0000000000000001",
	34177 => "0000000000000001",34178 => "0000000000000001",34179 => "0000000000000001",
	34180 => "0000000000000001",34181 => "0000000000000001",34182 => "0000000000000001",
	34183 => "0000000000000001",34184 => "0000000000000001",34185 => "0000000000000001",
	34186 => "0000000000000001",34187 => "0000000000000001",34188 => "0000000000000000",
	34189 => "0000000000000000",34190 => "0000000000000000",34191 => "0000000000000000",
	34192 => "0000000000000000",34193 => "0000000000000000",34194 => "0000000000000000",
	others =>"0000000000000000"
);

SIGNAL not_index,minus_index,zeros : std_logic_vector(15 downto 0);

begin
	
	zeros <= (others=>'0');

	not_index_map : for i in 0 to 15 GENERATE 
		not_map : not_index(i) <= not bitVector(i);
	end GENERATE;

	minus_index_map : fulladder_n 
		GENERIC MAP (n=>16)
		PORT MAP (
			cin => '1',
			x => not_index,
			y => zeros,
			z => minus_index
			);


	findValue: process (clk,bitVector) is 
		variable index : integer := 0;
		variable index_sign : integer := 0;
		variable temp_index : std_logic_vector(15 downto 0); 

		BEGIN  
			if bitVector(15)='1' then
				temp_index := '1'&minus_index(14 downto 0);
			else
				temp_index := bitVector;
			end if;

			index := to_integer(unsigned(temp_index));
			if index < 3000 then
				outVector <= exp_lut(index);
			else 
				if index > 32768 then
					--new_index := index - 32768;
					if index < 34190 then
						outVector <= exp_lut_neg(index);
					else
						outVector <= x"0000";
					end if;
				else 
					outVector <= x"0000";
				end if;
			end if;

	end process findValue;

end architecture;

